** sch_path: /foss/designs/libs/core_bandgap/bandgap/bandgap.sch
.subckt bandgap VDD VBG IPTAT IZTC SUB VSS vpref vpref_fb ICTAT VZTC
*.PININFO VDD:B VSS:B SUB:B VBG:B IPTAT:B IZTC:B vpref:B vpref_fb:B ICTAT:B VZTC:B
* noconn SUB
XQ1 VSS VSS vbe pnp_05p00x00p42 m=2
XQ2 VSS VSS vbjt_ptat[0] pnp_05p00x00p42 m=16
Mpref1 net2 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
Mpref2 net1 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
XRptat[5] vbjt_ptat[5] vbjt_ptat[6] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat[4] vbjt_ptat[4] vbjt_ptat[5] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat[3] vbjt_ptat[3] vbjt_ptat[4] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat[2] vbjt_ptat[2] vbjt_ptat[3] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat[1] vbjt_ptat[1] vbjt_ptat[2] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat[0] vbjt_ptat[0] vbjt_ptat[1] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
* tap: vbjt_ptat[5:0] --> vbjt_ptat[0]
* tap: vbjt_ptat[6:1] --> vbjt_ptat[6]
XQ3 VSS VSS vbjt_bg[0] pnp_05p00x00p42 m=2
Mpref3 net3 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
XRref[53] vbjt_bg[53] VBG VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[52] vbjt_bg[52] vbjt_bg[53] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[51] vbjt_bg[51] vbjt_bg[52] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[50] vbjt_bg[50] vbjt_bg[51] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[49] vbjt_bg[49] vbjt_bg[50] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[48] vbjt_bg[48] vbjt_bg[49] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[47] vbjt_bg[47] vbjt_bg[48] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[46] vbjt_bg[46] vbjt_bg[47] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[45] vbjt_bg[45] vbjt_bg[46] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[44] vbjt_bg[44] vbjt_bg[45] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[43] vbjt_bg[43] vbjt_bg[44] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[42] vbjt_bg[42] vbjt_bg[43] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[41] vbjt_bg[41] vbjt_bg[42] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[40] vbjt_bg[40] vbjt_bg[41] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[39] vbjt_bg[39] vbjt_bg[40] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[38] vbjt_bg[38] vbjt_bg[39] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[37] vbjt_bg[37] vbjt_bg[38] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[36] vbjt_bg[36] vbjt_bg[37] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[35] vbjt_bg[35] vbjt_bg[36] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[34] vbjt_bg[34] vbjt_bg[35] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[33] vbjt_bg[33] vbjt_bg[34] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[32] vbjt_bg[32] vbjt_bg[33] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[31] vbjt_bg[31] vbjt_bg[32] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[30] vbjt_bg[30] vbjt_bg[31] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[29] vbjt_bg[29] vbjt_bg[30] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[28] vbjt_bg[28] vbjt_bg[29] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[27] vbjt_bg[27] vbjt_bg[28] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[26] vbjt_bg[26] vbjt_bg[27] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[25] vbjt_bg[25] vbjt_bg[26] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[24] vbjt_bg[24] vbjt_bg[25] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[23] vbjt_bg[23] vbjt_bg[24] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[22] vbjt_bg[22] vbjt_bg[23] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[21] vbjt_bg[21] vbjt_bg[22] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[20] vbjt_bg[20] vbjt_bg[21] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[19] vbjt_bg[19] vbjt_bg[20] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[18] vbjt_bg[18] vbjt_bg[19] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[17] vbjt_bg[17] vbjt_bg[18] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[16] vbjt_bg[16] vbjt_bg[17] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[15] vbjt_bg[15] vbjt_bg[16] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[14] vbjt_bg[14] vbjt_bg[15] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[13] vbjt_bg[13] vbjt_bg[14] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[12] vbjt_bg[12] vbjt_bg[13] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[11] vbjt_bg[11] vbjt_bg[12] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[10] vbjt_bg[10] vbjt_bg[11] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[9] vbjt_bg[9] vbjt_bg[10] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[8] vbjt_bg[8] vbjt_bg[9] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[7] vbjt_bg[7] vbjt_bg[8] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[6] vbjt_bg[6] vbjt_bg[7] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[5] vbjt_bg[5] vbjt_bg[6] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[4] vbjt_bg[4] vbjt_bg[5] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[3] vbjt_bg[3] vbjt_bg[4] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[2] vbjt_bg[2] vbjt_bg[3] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[1] vbjt_bg[1] vbjt_bg[2] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRref[0] vbjt_bg[0] vbjt_bg[1] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
* tap: vbjt_bg[53:0] --> vbjt_bg[0]
Mpref4 net4 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
Mpref5 vbjt_ptat[6] vpcas net2 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
Mpref6 vbe vpcas net1 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
Mpref7 VBG vpcas net3 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
Mpref8 IPTAT vpcas net4 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
XQ4 VSS VSS vbe2 pnp_05p00x00p42 m=2
Mnref5 vnref_ctat vnref_ctat vbjt_ctat[34] vbjt_ctat[34] nfet_05v0 L=0.6u W=4u nf=1 m=16
Mnref6 vgs_ctat vnref_ctat vbe2 vbe2 nfet_05v0 L=0.6u W=4u nf=1 m=16
XRptat1[33] vbjt_ctat[33] vbjt_ctat[34] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[32] vbjt_ctat[32] vbjt_ctat[33] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[31] vbjt_ctat[31] vbjt_ctat[32] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[30] vbjt_ctat[30] vbjt_ctat[31] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[29] vbjt_ctat[29] vbjt_ctat[30] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[28] vbjt_ctat[28] vbjt_ctat[29] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[27] vbjt_ctat[27] vbjt_ctat[28] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[26] vbjt_ctat[26] vbjt_ctat[27] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[25] vbjt_ctat[25] vbjt_ctat[26] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[24] vbjt_ctat[24] vbjt_ctat[25] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[23] vbjt_ctat[23] vbjt_ctat[24] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[22] vbjt_ctat[22] vbjt_ctat[23] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[21] vbjt_ctat[21] vbjt_ctat[22] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[20] vbjt_ctat[20] vbjt_ctat[21] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[19] vbjt_ctat[19] vbjt_ctat[20] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[18] vbjt_ctat[18] vbjt_ctat[19] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[17] vbjt_ctat[17] vbjt_ctat[18] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[16] vbjt_ctat[16] vbjt_ctat[17] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[15] vbjt_ctat[15] vbjt_ctat[16] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[14] vbjt_ctat[14] vbjt_ctat[15] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[13] vbjt_ctat[13] vbjt_ctat[14] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[12] vbjt_ctat[12] vbjt_ctat[13] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[11] vbjt_ctat[11] vbjt_ctat[12] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[10] vbjt_ctat[10] vbjt_ctat[11] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[9] vbjt_ctat[9] vbjt_ctat[10] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[8] vbjt_ctat[8] vbjt_ctat[9] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[7] vbjt_ctat[7] vbjt_ctat[8] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[6] vbjt_ctat[6] vbjt_ctat[7] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[5] vbjt_ctat[5] vbjt_ctat[6] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[4] vbjt_ctat[4] vbjt_ctat[5] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[3] vbjt_ctat[3] vbjt_ctat[4] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[2] vbjt_ctat[2] vbjt_ctat[3] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[1] vbjt_ctat[1] vbjt_ctat[2] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat1[0] VSS vbjt_ctat[1] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
* tap: vbjt_ctat[34:1] --> vbjt_ctat[34]
Mnref7 vpcas_ctat vgs_ctat VSS VSS nfet_05v0 L=4u W=1u nf=1 m=1
Mpref9 net5 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
Mpref10 vgs_ctat vpcas net5 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
Mpref11 net6 vpref_ctat VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=4
Mpref12 net7 vpref_ctat VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=4
XRpcas1[7] vr_pcas_ctat[7] vpref_ctat VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[6] vr_pcas_ctat[6] vr_pcas_ctat[7] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[5] vr_pcas_ctat[5] vr_pcas_ctat[6] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[4] vr_pcas_ctat[4] vr_pcas_ctat[5] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[3] vr_pcas_ctat[3] vr_pcas_ctat[4] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[2] vr_pcas_ctat[2] vr_pcas_ctat[3] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[1] vr_pcas_ctat[1] vr_pcas_ctat[2] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRpcas1[0] vpcas_ctat vr_pcas_ctat[1] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
Mpref13 vpref_ctat vpcas_ctat net6 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=16
Mpref14 vnref_ctat vpcas_ctat net7 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=16
Mpref15 net8 vpref_ctat VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=6
Mpref16 VZTC vpcas_ctat net8 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=24
XRptat2[30] v_ztc[30] VZTC VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[29] v_ztc[29] v_ztc[30] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[28] v_ztc[28] v_ztc[29] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[27] v_ztc[27] v_ztc[28] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[26] v_ztc[26] v_ztc[27] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[25] v_ztc[25] v_ztc[26] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[24] v_ztc[24] v_ztc[25] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[23] v_ztc[23] v_ztc[24] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[22] v_ztc[22] v_ztc[23] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[21] v_ztc[21] v_ztc[22] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[20] v_ztc[20] v_ztc[21] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[19] v_ztc[19] v_ztc[20] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[18] v_ztc[18] v_ztc[19] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[17] v_ztc[17] v_ztc[18] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[16] v_ztc[16] v_ztc[17] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[15] v_ztc[15] v_ztc[16] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[14] v_ztc[14] v_ztc[15] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[13] v_ztc[13] v_ztc[14] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[12] v_ztc[12] v_ztc[13] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[11] v_ztc[11] v_ztc[12] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[10] v_ztc[10] v_ztc[11] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[9] v_ztc[9] v_ztc[10] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[8] v_ztc[8] v_ztc[9] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[7] v_ztc[7] v_ztc[8] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[6] v_ztc[6] v_ztc[7] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[5] v_ztc[5] v_ztc[6] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[4] v_ztc[4] v_ztc[5] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[3] v_ztc[3] v_ztc[4] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[2] v_ztc[2] v_ztc[3] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[1] v_ztc[1] v_ztc[2] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
XRptat2[0] VSS v_ztc[1] VDD ppolyf_u_1k r_width=1e-6 r_length=4.5e-6 m=1
Mpref17 net9 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
Mpref18 VZTC vpcas net9 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
Mpref_dumm_L[3] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_L[2] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_L[1] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_L[0] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_TP[17] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[16] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[15] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[14] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[13] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[12] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[11] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[10] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[9] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[8] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[7] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[6] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[5] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[4] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[3] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[2] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[1] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP[0] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
x1 VDD net12 vbe vbjt_ptat[6] vpref_fb VSS bandgap_opamp
Mpref19 net10 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
Mpref20 net11 vpcas net10 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
M1 net11 net11 VSS VSS nfet_05v0 L=2u W=0.5u nf=1 m=2
M2 net16 net11 VSS VSS nfet_05v0 L=2u W=0.5u nf=1 m=2
M3 vpcas net11 VSS VSS nfet_05v0 L=2u W=0.5u nf=1 m=2
Mpref21 vpcas vpcas VDD VDD pfet_05v0 L=3.2u W=3.2u nf=1 m=8
XRptat3[33] vbias[33] vstart_up VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[32] vbias[32] vbias[33] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[31] vbias[31] vbias[32] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[30] vbias[30] vbias[31] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[29] vbias[29] vbias[30] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[28] vbias[28] vbias[29] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[27] vbias[27] vbias[28] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[26] vbias[26] vbias[27] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[25] vbias[25] vbias[26] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[24] vbias[24] vbias[25] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[23] vbias[23] vbias[24] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[22] vbias[22] vbias[23] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[21] vbias[21] vbias[22] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[20] vbias[20] vbias[21] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[19] vbias[19] vbias[20] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[18] vbias[18] vbias[19] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[17] vbias[17] vbias[18] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[16] vbias[16] vbias[17] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[15] vbias[15] vbias[16] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[14] vbias[14] vbias[15] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[13] vbias[13] vbias[14] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[12] vbias[12] vbias[13] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[11] vbias[11] vbias[12] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[10] vbias[10] vbias[11] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[9] vbias[9] vbias[10] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[8] vbias[8] vbias[9] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[7] vbias[7] vbias[8] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[6] vbias[6] vbias[7] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[5] vbias[5] vbias[6] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[4] vbias[4] vbias[5] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[3] vbias[3] vbias[4] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[2] vbias[2] vbias[3] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[1] vbias[1] vbias[2] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
XRptat3[0] VSS vbias[1] VDD ppolyf_u_1k r_width=0.5e-6 r_length=4.5e-6 m=1
Mpref23 vstart_up vpcas VDD VDD pfet_05v0 L=0.5u W=4u nf=1 m=16
Mpref24 VSS vstart_up vpcas vpcas pfet_05v0 L=0.5u W=4u nf=1 m=32
Mpref25 net13 vpref_ctat VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=4
Mpref26 ICTAT vpcas_ctat net13 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=16
Mpref27 net14 vpref_ctat VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=6
Mpref28 IZTC vpcas_ctat net14 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=24
Mpref29 net15 vpref VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=2
Mpref30 IZTC vpcas net15 VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=8
M5 VSS vstart_up VSS VSS nfet_05v0 L=1u W=4u nf=1 m=32
M4 net12 vstart_up net16 VSS nfet_05v0 L=0.6u W=1u nf=1 m=1
Mpref22 VSS vstart_up vpref vpref pfet_05v0 L=0.5u W=4u nf=1 m=32
M6 VSS vgs_ctat VSS VSS nfet_05v0 L=1u W=3.2u nf=1 m=32
Mpcas_dumm_L[7] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[6] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[5] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[4] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[3] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[2] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[1] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L[0] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_TP[35] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[34] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[33] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[32] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[31] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[30] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[29] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[28] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[27] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[26] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[25] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[24] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[23] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[22] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[21] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[20] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[19] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[18] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[17] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[16] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[15] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[14] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[13] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[12] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[11] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[10] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[9] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[8] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[7] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[6] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[5] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[4] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[3] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[2] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[1] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP[0] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_L1[3] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_L1[2] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_L1[1] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_L1[0] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpref_dumm_TP1[19] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[18] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[17] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[16] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[15] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[14] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[13] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[12] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[11] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[10] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[9] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[8] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[7] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[6] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[5] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[4] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[3] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[2] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[1] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpref_dumm_TP1[0] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_L1[7] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[6] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[5] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[4] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[3] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[2] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[1] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_L1[0] VDD VDD VDD VDD pfet_05v0 L=0.8u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[39] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[38] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[37] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[36] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[35] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[34] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[33] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[32] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[31] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[30] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[29] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[28] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[27] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[26] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[25] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[24] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[23] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[22] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[21] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[20] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[19] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[18] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[17] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[16] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[15] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[14] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[13] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[12] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[11] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[10] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[9] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[8] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[7] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[6] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[5] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[4] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[3] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[2] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[1] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
Mpcas_dumm_TP1[0] VDD VDD VDD VDD pfet_05v0 L=0.6u W=3.2u nf=1 m=1
.ends

* expanding   symbol:  libs/core_bandgap/bandgap_opamp/bandgap_opamp.sym # of pins=6
** sym_path: /foss/designs/libs/core_bandgap/bandgap_opamp/bandgap_opamp.sym
** sch_path: /foss/designs/libs/core_bandgap/bandgap_opamp/bandgap_opamp.sch
.subckt bandgap_opamp VDD ibias vn vp vout VSS
*.PININFO vn:I vp:I vout:O ibias:I VDD:B VSS:B
Mpref0 ibias ibias VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=2
Mnload0 vnload vnload VSS VSS nfet_05v0 L=2u W=0.5u nf=1 m=2
Mpref1 vptail ibias VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=2
Mpref2 vout ibias VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=8
Mpdiff0 vnload vn vptail VDD pfet_05v0 L=1u W=2u nf=1 m=2
Mpdiff1 vout_1st vp vptail VDD pfet_05v0 L=1u W=2u nf=1 m=2
Mnload1 vout_1st vnload VSS VSS nfet_05v0 L=2u W=0.5u nf=1 m=2
Mncs vout vout_1st VSS VSS nfet_05v0 L=2u W=0.5u nf=1 m=16
Mpref_dumm_L[3] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_L[2] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_L[1] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_L[0] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[23] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[22] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[21] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[20] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[19] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[18] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[17] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[16] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[15] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[14] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[13] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[12] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[11] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[10] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[9] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[8] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[7] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[6] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[5] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[4] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[3] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[2] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[1] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
Mpref_dumm_TP[0] VDD VDD VDD VDD pfet_05v0 L=1u W=0.5u nf=1 m=1
XC1[5] vout vout_1st cap_mim_1f0fF c_width=10e-6 c_length=10e-6 m=1
XC1[4] vout vout_1st cap_mim_1f0fF c_width=10e-6 c_length=10e-6 m=1
XC1[3] vout vout_1st cap_mim_1f0fF c_width=10e-6 c_length=10e-6 m=1
XC1[2] vout vout_1st cap_mim_1f0fF c_width=10e-6 c_length=10e-6 m=1
XC1[1] vout vout_1st cap_mim_1f0fF c_width=10e-6 c_length=10e-6 m=1
XC1[0] vout vout_1st cap_mim_1f0fF c_width=10e-6 c_length=10e-6 m=1
.ends

