* Extracted by KLayout with GF180MCU LVS runset on : 21/08/2025 06:35

.SUBCKT bandgap I1_default_C I1_default_B I1_default_E SUB
M$1 \$386 \$433 \$385 \$456 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$2 \$388 \$434 \$387 \$454 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$3 \$390 \$435 \$389 \$452 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$4 \$392 \$436 \$391 \$450 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$5 \$394 \$437 \$393 \$447 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$6 \$396 \$438 \$395 \$445 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$7 \$398 \$439 \$397 \$444 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$8 \$400 \$440 \$399 \$442 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$9 \$466 \$529 \$465 \$551 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$10 \$468 \$530 \$467 \$547 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$11 \$470 \$531 \$469 \$544 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$12 \$472 \$532 \$471 \$542 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$13 \$474 \$533 \$473 \$560 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$14 \$476 \$534 \$475 \$557 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$15 \$478 \$535 \$477 \$555 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$16 \$480 \$536 \$479 \$553 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$17 \$562 \$601 \$561 \$622 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$18 \$564 \$602 \$563 \$626 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$19 \$566 \$603 \$565 \$631 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$20 \$568 \$604 \$567 \$624 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$21 \$570 \$605 \$569 \$676 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$22 \$572 \$606 \$571 \$673 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$23 \$574 \$607 \$573 \$672 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$24 \$576 \$608 \$575 \$670 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$25 \$686 \$781 \$685 \$823 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$26 \$688 \$782 \$687 \$822 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$27 \$690 \$783 \$689 \$819 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$28 \$692 \$784 \$691 \$818 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$29 \$694 \$785 \$693 \$815 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$30 \$696 \$786 \$695 \$814 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$31 \$698 \$787 \$697 \$812 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$32 \$700 \$788 \$699 \$809 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$33 \$850 \$893 \$849 \$940 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$34 \$852 \$894 \$851 \$945 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$35 \$854 \$895 \$853 \$946 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$36 \$856 \$896 \$855 \$951 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$37 \$858 \$897 \$857 \$952 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$38 \$860 \$898 \$859 \$957 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$39 \$862 \$899 \$861 \$958 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$40 \$864 \$900 \$863 \$937 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$41 \$1006 \$1067 \$1005 \$1075 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$42 \$1008 \$1068 \$1007 \$1079 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$43 \$1010 \$1069 \$1009 \$1082 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$44 \$1012 \$1070 \$1011 \$1085 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$45 \$1014 \$1071 \$1013 \$1126 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$46 \$1016 \$1072 \$1015 \$1128 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$47 \$1018 \$1073 \$1017 \$1130 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$48 \$1020 \$1074 \$1019 \$1132 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$49 \$1154 \$1290 \$1153 \$1308 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$50 \$1156 \$1291 \$1155 \$1310 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$51 \$1158 \$1292 \$1157 \$1314 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$52 \$1160 \$1293 \$1159 \$1316 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$53 \$1162 \$1294 \$1161 \$1320 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$54 \$1164 \$1295 \$1163 \$1322 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$55 \$1166 \$1296 \$1165 \$1325 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$56 \$1168 \$1297 \$1167 \$1328 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$57 \$1379 \$1450 \$1378 \$1477 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$58 \$1381 \$1451 \$1380 \$1480 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$59 \$1383 \$1452 \$1382 \$1473 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$60 \$1385 \$1453 \$1384 \$1470 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$61 \$1387 \$1454 \$1386 \$1467 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$62 \$1389 \$1455 \$1388 \$1464 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$63 \$1391 \$1456 \$1390 \$1462 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$64 \$1393 \$1457 \$1392 \$1459 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$65 \$1518 \$1618 \$1517 \$1651 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$66 \$1520 \$1619 \$1519 \$1654 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$67 \$1522 \$1620 \$1521 \$1658 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$68 \$1524 \$1621 \$1523 \$1664 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$69 \$1526 \$1622 \$1525 \$1667 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$70 \$1528 \$1623 \$1527 \$1669 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$71 \$1530 \$1624 \$1529 \$1675 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$72 \$1532 \$1625 \$1531 \$1677 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$73 \$1534 \$1626 \$1533 \$1681 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$74 \$1536 \$1627 \$1535 \$1684 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$75 \$1559 \$1628 \$1558 \$1687 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$76 \$1561 \$1629 \$1560 \$1692 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$77 \$1563 \$1630 \$1562 \$1694 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$78 \$1565 \$1631 \$1564 \$1697 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$79 \$1567 \$1632 \$1566 \$1701 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$80 \$1569 \$1633 \$1568 \$1704 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$81 \$1571 \$1634 \$1570 \$1706 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$82 \$1573 \$1635 \$1572 \$1710 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$83 \$1575 \$1636 \$1574 \$1712 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$84 \$1577 \$1637 \$1576 \$1715 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$85 \$1579 \$1638 \$1578 \$1718 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$86 \$1581 \$1639 \$1580 \$1722 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$87 \$1583 \$1640 \$1582 \$1724 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$88 \$1585 \$1641 \$1584 \$1727 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$89 \$1587 \$1642 \$1586 \$1672 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$90 \$1589 \$1643 \$1588 \$1662 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$91 \$1730 \$1836 \$1729 \$1872 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$92 \$1732 \$1837 \$1731 \$1873 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$93 \$1734 \$1838 \$1733 \$1876 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$94 \$1736 \$1839 \$1735 \$1881 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$95 \$1738 \$1840 \$1737 \$1888 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$96 \$1740 \$1841 \$1739 \$1892 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$97 \$1742 \$1842 \$1741 \$1897 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$98 \$1744 \$1843 \$1743 \$1901 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$99 \$1746 \$1844 \$1745 \$1906 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$100 \$1748 \$1845 \$1747 \$1909 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$101 \$1750 \$1846 \$1749 \$1916 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$102 \$1752 \$1847 \$1751 \$1922 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$103 \$1754 \$1848 \$1753 \$1923 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$104 \$1756 \$1849 \$1755 \$1928 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$105 \$1758 \$1850 \$1757 \$1930 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$106 \$1760 \$1851 \$1759 \$1934 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$107 \$1762 \$1852 \$1761 \$1936 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$108 \$1764 \$1853 \$1763 \$1940 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$109 \$1766 \$1854 \$1765 \$1943 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$110 \$1768 \$1855 \$1767 \$1946 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$111 \$1770 \$1856 \$1769 \$1949 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$112 \$1772 \$1857 \$1771 \$1952 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$113 \$1774 \$1858 \$1773 \$1919 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$114 \$1776 \$1859 \$1775 \$1912 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$115 \$1778 \$1860 \$1777 \$1902 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$116 \$1780 \$1861 \$1779 \$1893 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$117 \$1782 \$1862 \$1781 \$1884 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$118 \$1784 \$1863 \$1783 \$1883 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$119 \$2027 \$2068 \$2026 \$2104 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$120 \$2029 \$2069 \$2028 \$2108 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$121 \$1954 \$2070 \$1953 \$2109 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$122 \$1956 \$2071 \$1955 \$2115 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$123 \$1958 \$2072 \$1957 \$2120 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$124 \$1960 \$2073 \$1959 \$2122 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$125 \$1962 \$2074 \$1961 \$2127 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$126 \$1964 \$2075 \$1963 \$2132 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$127 \$1966 \$2076 \$1965 \$2134 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$128 \$1968 \$2077 \$1967 \$2138 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$129 \$1970 \$2078 \$1969 \$2141 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$130 \$1972 \$2079 \$1971 \$2145 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$131 \$1974 \$2080 \$1973 \$2150 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$132 \$1976 \$2081 \$1975 \$2153 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$133 \$1978 \$2082 \$1977 \$2157 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$134 \$1980 \$2083 \$1979 \$2159 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$135 \$1982 \$2084 \$1981 \$2163 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$136 \$1984 \$2085 \$1983 \$2166 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$137 \$1986 \$2086 \$1985 \$2168 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$138 \$1988 \$2087 \$1987 \$2172 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$139 \$1990 \$2088 \$1989 \$2175 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$140 \$1992 \$2089 \$1991 \$2148 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$141 \$1994 \$2090 \$1993 \$2142 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$142 \$1996 \$2091 \$1995 \$2136 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$143 \$1998 \$2092 \$1997 \$2129 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$144 \$2000 \$2093 \$1999 \$2123 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$145 \$2002 \$2094 \$2001 \$2117 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$146 \$2004 \$2095 \$2003 \$2112 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$147 \$2289 \$2395 \$2288 \$2465 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$148 \$2291 \$2396 \$2290 \$2467 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$149 \$2178 \$2292 \$2177 \$2329 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$150 \$2180 \$2293 \$2179 \$2332 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$151 \$2182 \$2294 \$2181 \$2334 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$152 \$2184 \$2295 \$2183 \$2335 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$153 \$2186 \$2296 \$2185 \$2337 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$154 \$2188 \$2297 \$2187 \$2340 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$155 \$2190 \$2298 \$2189 \$2342 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$156 \$2192 \$2299 \$2191 \$2343 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$157 \$2194 \$2300 \$2193 \$2346 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$158 \$2196 \$2301 \$2195 \$2347 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$159 \$2198 \$2302 \$2197 \$2352 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$160 \$2200 \$2303 \$2199 \$2355 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$161 \$2202 \$2304 \$2201 \$2361 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$162 \$2204 \$2305 \$2203 \$2366 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$163 \$2206 \$2306 \$2205 \$2370 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$164 \$2208 \$2307 \$2207 \$2372 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$165 \$2210 \$2308 \$2209 \$2379 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$166 \$2212 \$2309 \$2211 \$2383 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$167 \$2214 \$2310 \$2213 \$2387 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$168 \$2216 \$2311 \$2215 \$2390 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$169 \$2218 \$2312 \$2217 \$2392 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$170 \$2220 \$2313 \$2219 \$2384 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$171 \$2222 \$2314 \$2221 \$2375 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$172 \$2224 \$2315 \$2223 \$2363 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$173 \$2226 \$2316 \$2225 \$2354 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$174 \$2228 \$2317 \$2227 \$2328 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$175 \$2451 \$2626 \$2450 \$2663 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$176 \$2453 \$2627 \$2452 \$2665 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$177 \$2455 \$2628 \$2454 \$2666 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$178 \$2457 \$2629 \$2456 \$2668 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$179 \$2398 \$2490 \$2397 \$2529 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$180 \$2400 \$2491 \$2399 \$2533 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$181 \$2402 \$2492 \$2401 \$2536 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$182 \$2404 \$2493 \$2403 \$2538 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$183 \$2406 \$2494 \$2405 \$2542 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$184 \$2408 \$2495 \$2407 \$2545 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$185 \$2410 \$2496 \$2409 \$2548 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$186 \$2412 \$2497 \$2411 \$2551 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$187 \$2414 \$2498 \$2413 \$2553 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$188 \$2416 \$2499 \$2415 \$2557 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$189 \$2418 \$2500 \$2417 \$2559 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$190 \$2420 \$2501 \$2419 \$2526 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$191 \$2422 \$2502 \$2421 \$2522 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$192 \$2424 \$2503 \$2423 \$2520 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$193 \$2426 \$2504 \$2425 \$2516 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$194 \$2428 \$2505 \$2427 \$2515 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$195 \$2562 \$2691 \$2561 \$2725 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$196 \$2564 \$2692 \$2563 \$2728 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$197 \$2566 \$2693 \$2565 \$2731 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$198 \$2568 \$2694 \$2567 \$2734 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$199 \$2570 \$2695 \$2569 \$2736 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$200 \$2572 \$2696 \$2571 \$2739 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$201 \$2574 \$2697 \$2573 \$2742 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$202 \$2576 \$2698 \$2575 \$2746 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$203 \$2578 \$2699 \$2577 \$2749 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$204 \$2580 \$2700 \$2579 \$2752 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$205 \$2582 \$2701 \$2581 \$2754 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$206 \$2584 \$2702 \$2583 \$2758 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$207 \$2586 \$2703 \$2585 \$2760 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$208 \$2588 \$2704 \$2587 \$2764 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$209 \$2590 \$2705 \$2589 \$2767 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$210 \$2592 \$2706 \$2591 \$2769 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$211 \$2594 \$2707 \$2593 \$2773 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$212 \$2596 \$2708 \$2595 \$2775 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$213 \$2598 \$2709 \$2597 \$2779 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$214 \$2600 \$2710 \$2599 \$2781 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$215 \$2795 \$2950 \$2794 \$3006 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$216 \$2797 \$2951 \$2796 \$3009 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$217 \$2799 \$2952 \$2798 \$3011 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$218 \$2801 \$2953 \$2800 \$3012 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$219 \$2858 \$2954 \$2857 \$3018 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$220 \$2860 \$2955 \$2859 \$3021 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$221 \$2862 \$2956 \$2861 \$3025 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$222 \$2864 \$2957 \$2863 \$3027 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$223 \$2866 \$2958 \$2865 \$3030 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$224 \$2868 \$2959 \$2867 \$3033 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$225 \$2870 \$2960 \$2869 \$3036 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$226 \$2872 \$2961 \$2871 \$3039 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$227 \$2874 \$2962 \$2873 \$3042 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$228 \$2876 \$2963 \$2875 \$3045 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$229 \$2878 \$2964 \$2877 \$3048 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$230 \$2880 \$2965 \$2879 \$3015 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$231 \$2882 \$2966 \$2881 \$3003 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$232 \$2884 \$2967 \$2883 \$3000 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$233 \$2886 \$2968 \$2885 \$2997 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$234 \$2888 \$2969 \$2887 \$2995 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$235 \$2890 \$2970 \$2889 \$2992 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$236 \$2892 \$2971 \$2891 \$2989 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$237 \$2631 \$2802 \$2630 \$2856 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$238 \$2633 \$2803 \$2632 \$2853 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$239 \$2635 \$2804 \$2634 \$2852 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$240 \$2637 \$2805 \$2636 \$2850 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$241 \$2639 \$2806 \$2638 \$2847 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$242 \$2641 \$2807 \$2640 \$2845 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$243 \$2643 \$2808 \$2642 \$2844 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$244 \$2645 \$2809 \$2644 \$2841 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$245 \$2647 \$2810 \$2646 \$2839 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$246 \$2649 \$2811 \$2648 \$2837 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$247 \$2651 \$2812 \$2650 \$2836 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$248 \$2653 \$2813 \$2652 \$2834 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$249 \$2655 \$2814 \$2654 \$2831 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$250 \$2657 \$2815 \$2656 \$2830 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$251 \$2659 \$2816 \$2658 \$2827 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$252 \$2661 \$2817 \$2660 \$2825 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$253 \$2915 \$3050 \$2914 \$3060 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$254 \$2917 \$3051 \$2916 \$3062 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$255 \$3074 \$3130 \$3073 \$3260 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$256 \$3076 \$3131 \$3075 \$3257 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$257 \$3078 \$3132 \$3077 \$3256 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$258 \$3080 \$3133 \$3079 \$3254 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$259 \$3082 \$3134 \$3081 \$3251 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$260 \$3084 \$3135 \$3083 \$3249 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$261 \$3086 \$3136 \$3085 \$3248 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$262 \$3088 \$3137 \$3087 \$3245 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$263 \$3090 \$3138 \$3089 \$3243 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$264 \$3092 \$3139 \$3091 \$3242 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$265 \$3094 \$3140 \$3093 \$3240 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$266 \$3096 \$3141 \$3095 \$3238 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$267 \$3098 \$3142 \$3097 \$3235 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$268 \$3100 \$3143 \$3099 \$3233 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$269 \$3102 \$3144 \$3101 \$3232 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$270 \$3104 \$3145 \$3103 \$3230 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$271 \$3106 \$3146 \$3105 \$3227 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$272 \$3108 \$3147 \$3107 \$3226 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$273 \$2973 \$3148 \$2972 \$3193 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$274 \$2975 \$3149 \$2974 \$3187 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$275 \$2977 \$3150 \$2976 \$3182 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$276 \$2979 \$3151 \$2978 \$3178 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$277 \$2981 \$3152 \$2980 \$3173 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$278 \$2983 \$3153 \$2982 \$3170 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$279 \$2985 \$3154 \$2984 \$3167 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$280 \$2987 \$3155 \$2986 \$3163 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$281 \$3066 \$3282 \$3065 \$3295 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$282 \$3068 \$3283 \$3067 \$3296 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$283 \$3070 \$3284 \$3069 \$3300 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$284 \$3072 \$3285 \$3071 \$3303 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$285 \$3206 \$3372 \$3205 \$3419 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$286 \$3208 \$3373 \$3207 \$3421 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$287 \$3306 \$3374 \$3305 \$3502 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$288 \$3308 \$3375 \$3307 \$3504 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$289 \$3310 \$3376 \$3309 \$3499 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$290 \$3312 \$3377 \$3311 \$3497 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$291 \$3314 \$3378 \$3313 \$3495 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$292 \$3316 \$3379 \$3315 \$3493 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$293 \$3318 \$3380 \$3317 \$3492 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$294 \$3320 \$3381 \$3319 \$3489 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$295 \$3322 \$3382 \$3321 \$3487 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$296 \$3324 \$3383 \$3323 \$3486 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$297 \$3326 \$3384 \$3325 \$3484 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$298 \$3328 \$3385 \$3327 \$3481 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$299 \$3330 \$3386 \$3329 \$3480 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$300 \$3332 \$3387 \$3331 \$3478 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$301 \$3334 \$3388 \$3333 \$3476 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$302 \$3336 \$3389 \$3335 \$3474 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$303 \$3338 \$3390 \$3337 \$3471 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$304 \$3340 \$3391 \$3339 \$3470 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$305 \$3210 \$3392 \$3209 \$3438 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$306 \$3212 \$3393 \$3211 \$3434 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$307 \$3214 \$3394 \$3213 \$3429 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$308 \$3216 \$3395 \$3215 \$3425 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$309 \$3218 \$3396 \$3217 \$3416 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$310 \$3220 \$3397 \$3219 \$3413 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$311 \$3222 \$3398 \$3221 \$3412 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$312 \$3224 \$3399 \$3223 \$3407 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$313 \$3365 \$3594 \$3364 \$3614 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$314 \$3367 \$3595 \$3366 \$3616 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$315 \$3369 \$3596 \$3368 \$3621 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$316 \$3371 \$3597 \$3370 \$3623 pfet_05v0 L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$317 \$3534 \$3649 \$3533 \$3681 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$318 \$3536 \$3650 \$3535 \$3684 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$319 \$3538 \$3651 \$3537 \$3688 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$320 \$3540 \$3652 \$3539 \$3691 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$321 \$3542 \$3653 \$3541 \$3695 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$322 \$3544 \$3654 \$3543 \$3697 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$323 \$3546 \$3655 \$3545 \$3701 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$324 \$3548 \$3656 \$3547 \$3703 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$325 \$3550 \$3657 \$3549 \$3706 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$326 \$3552 \$3658 \$3551 \$3710 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$327 \$3554 \$3659 \$3553 \$3712 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$328 \$3556 \$3660 \$3555 \$3715 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$329 \$3558 \$3661 \$3557 \$3719 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$330 \$3560 \$3662 \$3559 \$3721 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$331 \$3562 \$3663 \$3561 \$3725 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$332 \$3564 \$3664 \$3563 \$3727 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$333 \$3566 \$3665 \$3565 \$3678 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$334 \$3568 \$3666 \$3567 \$3675 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$335 \$3570 \$3667 \$3569 \$3672 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$336 \$3572 \$3668 \$3571 \$3670 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$337 \$3454 \$3598 \$3453 \$3648 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$338 \$3456 \$3599 \$3455 \$3643 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$339 \$3458 \$3600 \$3457 \$3640 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$340 \$3460 \$3601 \$3459 \$3637 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$341 \$3462 \$3602 \$3461 \$3635 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$342 \$3464 \$3603 \$3463 \$3631 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$343 \$3466 \$3604 \$3465 \$3629 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$344 \$3468 \$3605 \$3467 \$3626 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$345 \$3839 \$3961 \$3838 \$3964 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$346 \$3841 \$3962 \$3840 \$3966 pfet_05v0 L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$347 \$3795 \$3842 \$3794 \$3898 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$348 \$3797 \$3843 \$3796 \$3901 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$349 \$3799 \$3844 \$3798 \$3905 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$350 \$3801 \$3845 \$3800 \$3907 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$351 \$3803 \$3846 \$3802 \$3911 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$352 \$3805 \$3847 \$3804 \$3913 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$353 \$3807 \$3848 \$3806 \$3916 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$354 \$3809 \$3849 \$3808 \$3919 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$355 \$3811 \$3850 \$3810 \$3923 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$356 \$3813 \$3851 \$3812 \$3925 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$357 \$3815 \$3852 \$3814 \$3928 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$358 \$3817 \$3853 \$3816 \$3932 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$359 \$3819 \$3854 \$3818 \$3934 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$360 \$3821 \$3855 \$3820 \$3938 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$361 \$3823 \$3856 \$3822 \$3941 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$362 \$3825 \$3857 \$3824 \$3943 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$363 \$3827 \$3858 \$3826 \$3946 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$364 \$3829 \$3859 \$3828 \$3949 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$365 \$3862 \$3969 \$3860 \$3979 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$366 \$3751 \$3861 \$3750 \$3952 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$367 \$3865 \$3970 \$3863 \$3985 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$368 \$3753 \$3864 \$3752 \$3958 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$369 \$3868 \$3971 \$3866 \$3991 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$370 \$3755 \$3867 \$3754 \$3959 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$371 \$3757 \$3870 \$3756 \$3956 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$372 \$3871 \$3972 \$3869 \$3995 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$373 \$3874 \$3973 \$3872 \$4000 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$374 \$3759 \$3873 \$3758 \$3953 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$375 \$3877 \$3974 \$3875 \$3994 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$376 \$3761 \$3876 \$3760 \$3895 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$377 \$3880 \$3975 \$3878 \$3987 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$378 \$3763 \$3879 \$3762 \$3893 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$379 \$3765 \$3882 \$3764 \$3891 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$380 \$3883 \$3976 \$3881 \$3980 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$381 \$4002 \$4017 \$4001 \$4027 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$382 \$4004 \$4018 \$4003 \$4030 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$383 \$4006 \$4019 \$4005 \$4033 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$384 \$4008 \$4020 \$4007 \$4035 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$385 \$4010 \$4021 \$4009 \$4039 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$386 \$4012 \$4022 \$4011 \$4042 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$387 \$4014 \$4023 \$4013 \$4044 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$388 \$4016 \$4024 \$4015 \$4047 pfet_05v0 L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$389 \$2 \$33 \$1 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$390 \$4 \$34 \$3 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$391 \$6 \$35 \$5 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$392 \$8 \$36 \$7 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$393 \$10 \$37 \$9 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$394 \$12 \$38 \$11 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$395 \$14 \$39 \$13 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$396 \$16 \$40 \$15 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$397 \$18 \$73 \$17 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$398 \$20 \$74 \$19 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$399 \$22 \$75 \$21 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$400 \$24 \$76 \$23 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$401 \$26 \$77 \$25 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$402 \$28 \$78 \$27 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$403 \$30 \$79 \$29 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$404 \$32 \$80 \$31 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$405 \$58 \$97 \$57 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$406 \$60 \$98 \$59 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$407 \$62 \$99 \$61 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U PD=9.46U
M$408 \$64 \$100 \$63 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$409 \$66 \$101 \$65 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$410 \$68 \$102 \$67 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$411 \$70 \$103 \$69 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$412 \$72 \$104 \$71 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$413 \$82 \$105 \$81 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$414 \$84 \$106 \$83 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$415 \$86 \$107 \$85 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$416 \$88 \$108 \$87 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$417 \$90 \$109 \$89 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$418 \$92 \$110 \$91 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$419 \$94 \$111 \$93 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$420 \$96 \$112 \$95 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$421 \$146 \$201 \$145 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$422 \$148 \$202 \$147 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$423 \$150 \$203 \$149 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$424 \$152 \$204 \$151 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$425 \$154 \$205 \$153 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$426 \$156 \$206 \$155 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$427 \$158 \$207 \$157 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$428 \$160 \$208 \$159 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$429 \$186 \$241 \$185 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$430 \$188 \$242 \$187 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$431 \$190 \$243 \$189 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$432 \$192 \$244 \$191 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$433 \$194 \$245 \$193 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$434 \$196 \$246 \$195 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$435 \$198 \$247 \$197 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$436 \$200 \$248 \$199 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$437 \$226 \$297 \$225 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$438 \$228 \$298 \$227 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$439 \$230 \$299 \$229 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$440 \$232 \$300 \$231 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$441 \$234 \$301 \$233 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$442 \$236 \$302 \$235 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$443 \$238 \$303 \$237 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$444 \$240 \$304 \$239 SUB nfet_05v0 L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$445 \$258 \$337 \$257 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$446 \$260 \$338 \$259 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$447 \$262 \$339 \$261 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$448 \$264 \$340 \$263 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$449 \$266 \$341 \$265 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$450 \$268 \$342 \$267 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$451 \$270 \$343 \$269 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$452 \$272 \$344 \$271 SUB nfet_05v0 L=1U W=3.2U AS=2.336P AD=2.336P PS=7.86U
+ PD=7.86U
M$453 \$722 \$789 \$721 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$454 \$634 \$701 \$633 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$455 \$724 \$790 \$723 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$456 \$636 \$702 \$635 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$457 \$638 \$703 \$637 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$458 \$726 \$791 \$725 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$459 \$640 \$704 \$639 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$460 \$728 \$792 \$727 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$461 \$642 \$705 \$641 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$462 \$730 \$793 \$729 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$463 \$644 \$706 \$643 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$464 \$732 \$794 \$731 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$465 \$646 \$707 \$645 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$466 \$734 \$795 \$733 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$467 \$736 \$796 \$735 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$468 \$648 \$708 \$647 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$469 \$738 \$797 \$737 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$470 \$650 \$709 \$649 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$471 \$740 \$798 \$739 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$472 \$652 \$710 \$651 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$473 \$866 \$905 \$865 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$474 \$868 \$906 \$867 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$475 \$870 \$907 \$869 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$476 \$872 \$908 \$871 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$477 \$874 \$909 \$873 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$478 \$876 \$910 \$875 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$479 \$878 \$911 \$877 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$480 \$880 \$912 \$879 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$481 \$882 \$913 \$881 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$482 \$884 \$914 \$883 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$483 \$886 \$901 \$885 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$484 \$888 \$902 \$887 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$485 \$890 \$903 \$889 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$486 \$892 \$904 \$891 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$487 \$982 \$1042 \$981 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$488 \$984 \$1043 \$983 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$489 \$986 \$1044 \$985 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$490 \$988 \$1045 \$987 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$491 \$990 \$1046 \$989 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$492 \$992 \$1047 \$991 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$493 \$994 \$1048 \$993 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$494 \$996 \$1049 \$995 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$495 \$998 \$1050 \$997 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$496 \$1000 \$1051 \$999 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$497 \$1025 \$1024 \$1023 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$498 \$971 \$970 \$969 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$499 \$1028 \$1027 \$1026 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$500 \$974 \$973 \$972 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$501 \$1031 \$1030 \$1029 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$502 \$977 \$976 \$975 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$503 \$1034 \$1033 \$1032 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$504 \$980 \$979 \$978 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$505 \$1022 \$1041 \$1021 SUB nfet_05v0 L=4U W=1U AS=0.73P AD=0.73P PS=3.46U
+ PD=3.46U
M$506 \$1106 \$1179 \$1105 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$507 \$1108 \$1180 \$1107 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$508 \$1110 \$1181 \$1109 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$509 \$1112 \$1182 \$1111 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$510 \$1114 \$1183 \$1113 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$511 \$1116 \$1184 \$1115 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$512 \$1118 \$1185 \$1117 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$513 \$1120 \$1186 \$1119 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$514 \$1122 \$1187 \$1121 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$515 \$1124 \$1188 \$1123 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$516 \$1146 \$1169 \$1145 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$517 \$1095 \$1094 \$1093 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$518 \$1148 \$1170 \$1147 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$519 \$1098 \$1097 \$1096 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$520 \$1101 \$1100 \$1099 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$521 \$1150 \$1171 \$1149 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$522 \$1104 \$1103 \$1102 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$523 \$1152 \$1172 \$1151 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$524 \$1239 \$1330 \$1238 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$525 \$1241 \$1331 \$1240 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$526 \$1243 \$1332 \$1242 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$527 \$1245 \$1333 \$1244 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$528 \$1247 \$1334 \$1246 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$529 \$1249 \$1335 \$1248 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$530 \$1251 \$1336 \$1250 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$531 \$1253 \$1337 \$1252 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$532 \$1255 \$1338 \$1254 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$533 \$1257 \$1339 \$1256 SUB nfet_05v0 L=0.6U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$534 \$1228 \$1227 \$1226 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$535 \$1231 \$1230 \$1229 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$536 \$1234 \$1233 \$1232 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$537 \$1237 \$1236 \$1235 SUB nfet_05v0 L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
Q$538 I1_default_C I1_default_B I1_default_E pnp_05p00x05p00 AE=1200P PE=960U
+ AB=41.9904P PB=25.92U AC=41.9904P PC=25.92U NE=48
R$586 \$1036 \$1037 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$587 \$1039 \$1040 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$588 \$1138 \$1139 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$589 \$1141 \$1142 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$590 \$1174 \$1175 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$591 \$1177 \$1178 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$592 \$1299 \$1300 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$593 \$1302 \$1303 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$594 \$1204 \$1205 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$595 \$1207 \$1208 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$596 \$1210 \$1211 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$597 \$1213 \$1214 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$598 \$1216 \$1217 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$599 \$1219 \$1220 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$600 \$1222 \$1223 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$601 \$1270 \$1271 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$602 \$1273 \$1274 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$603 \$1276 \$1277 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$604 \$1279 \$1280 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$605 \$1282 \$1283 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$606 \$1285 \$1286 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$607 \$1288 \$1289 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$608 \$1358 \$1359 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$609 \$1402 \$1403 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$610 \$1361 \$1362 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$611 \$1405 \$1406 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$612 \$1364 \$1365 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$613 \$1408 \$1409 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$614 \$1367 \$1368 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$615 \$1411 \$1412 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$616 \$1370 \$1371 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$617 \$1414 \$1415 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$618 \$1417 \$1418 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$619 \$1373 \$1374 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$620 \$1420 \$1421 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$621 \$1376 \$1377 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$622 \$1490 \$1491 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$623 \$1430 \$1431 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$624 \$1493 \$1494 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$625 \$1433 \$1434 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$626 \$1436 \$1437 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$627 \$1496 \$1497 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$628 \$1439 \$1440 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$629 \$1499 \$1500 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$630 \$1442 \$1443 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$631 \$1502 \$1503 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$632 \$1445 \$1446 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$633 \$1505 \$1506 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$634 \$1448 \$1449 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$635 \$1508 \$1509 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$636 \$1538 \$1539 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$637 \$1598 \$1599 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$638 \$1541 \$1542 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$639 \$1601 \$1602 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$640 \$1604 \$1605 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$641 \$1544 \$1545 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$642 \$1547 \$1548 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$643 \$1607 \$1608 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$644 \$1610 \$1611 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$645 \$1550 \$1551 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$646 \$1613 \$1614 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$647 \$1553 \$1554 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$648 \$1556 \$1557 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$649 \$1616 \$1617 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$650 \$1786 \$1787 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$651 \$1789 \$1790 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$652 \$1792 \$1793 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$653 \$1795 \$1796 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$654 \$1798 \$1799 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$655 \$1801 \$1802 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$656 \$1804 \$1805 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$657 \$1816 \$1817 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$658 \$2006 \$2007 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$659 \$2009 \$2010 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$660 \$1819 \$1820 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$661 \$2012 \$2013 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$662 \$1822 \$1823 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$663 \$2015 \$2016 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$664 \$1825 \$1826 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$665 \$1828 \$1829 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$666 \$2018 \$2019 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$667 \$2021 \$2022 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$668 \$1831 \$1832 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$669 \$1834 \$1835 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$670 \$2024 \$2025 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$671 \$2048 \$2049 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$672 \$2051 \$2052 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$673 \$2054 \$2055 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$674 \$2057 \$2058 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$675 \$2060 \$2061 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$676 \$2063 \$2064 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$677 \$2066 \$2067 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$678 \$2230 \$2231 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$679 \$2268 \$2269 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$680 \$2233 \$2234 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$681 \$2271 \$2272 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$682 \$2274 \$2275 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$683 \$2236 \$2237 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$684 \$2277 \$2278 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$685 \$2239 \$2240 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$686 \$2280 \$2281 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$687 \$2242 \$2243 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$688 \$2245 \$2246 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$689 \$2283 \$2284 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$690 \$2248 \$2249 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$691 \$2286 \$2287 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$692 \$2430 \$2431 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$693 \$2470 \$2471 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$694 \$2473 \$2474 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$695 \$2433 \$2434 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$696 \$2476 \$2477 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$697 \$2436 \$2437 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$698 \$2439 \$2440 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$699 \$2479 \$2480 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$700 \$2442 \$2443 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$701 \$2482 \$2483 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$702 \$2485 \$2486 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$703 \$2445 \$2446 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$704 \$2448 \$2449 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$705 \$2488 \$2489 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$706 \$2606 \$2607 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$707 \$2609 \$2610 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$708 \$2612 \$2613 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$709 \$2615 \$2616 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$710 \$2618 \$2619 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$711 \$2621 \$2622 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$712 \$2624 \$2625 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$713 \$2894 \$2895 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$714 \$2671 \$2672 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$715 \$2897 \$2898 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$716 \$2674 \$2675 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$717 \$2677 \$2678 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$718 \$2900 \$2901 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$719 \$2903 \$2904 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$720 \$2680 \$2681 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$721 \$2906 \$2907 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$722 \$2683 \$2684 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$723 \$2909 \$2910 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$724 \$2686 \$2687 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$725 \$2912 \$2913 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$726 \$2689 \$2690 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$727 \$2930 \$2931 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$728 \$2933 \$2934 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$729 \$2936 \$2937 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$730 \$2939 \$2940 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$731 \$2942 \$2943 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$732 \$2945 \$2946 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$733 \$2948 \$2949 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$734 \$3110 \$3111 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$735 \$3113 \$3114 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$736 \$3116 \$3117 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$737 \$3119 \$3120 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$738 \$3122 \$3123 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$739 \$3125 \$3126 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$740 \$3128 \$3129 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$741 \$3262 \$3263 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$742 \$3265 \$3266 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$743 \$3268 \$3269 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$744 \$3271 \$3272 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$745 \$3274 \$3275 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$746 \$3277 \$3278 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$747 \$3280 \$3281 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$748 \$3344 \$3345 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$749 \$3347 \$3348 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$750 \$3350 \$3351 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$751 \$3353 \$3354 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$752 \$3356 \$3357 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$753 \$3359 \$3360 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$754 \$3362 \$3363 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$755 \$3506 \$3507 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$756 \$3509 \$3510 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$757 \$3512 \$3513 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$758 \$3515 \$3516 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$759 \$3518 \$3519 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$760 \$3521 \$3522 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$761 \$3524 \$3525 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$762 \$3574 \$3575 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$763 \$3730 \$3731 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$764 \$3733 \$3734 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$765 \$3577 \$3578 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$766 \$3580 \$3581 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$767 \$3736 \$3737 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$768 \$3583 \$3584 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$769 \$3739 \$3740 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$770 \$3586 \$3587 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$771 \$3742 \$3743 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$772 \$3589 \$3590 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$773 \$3745 \$3746 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$774 \$3748 \$3749 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$775 \$3592 \$3593 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$776 \$3774 \$3775 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$777 \$3777 \$3778 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$778 \$3780 \$3781 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$779 \$3783 \$3784 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$780 \$3786 \$3787 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$781 \$3789 \$3790 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
R$782 \$3792 \$3793 SUB 4500 ppolyf_u_1k_6p0 L=4.5U W=1U
.ENDS bandgap
