** sch_path: /foss/designs/libs/core_top/top_amux_2x1/top_amux_2x1.sch
.subckt top_amux_2x1 IN0 VDD OUT VSS IN1 EN
*.PININFO VDD:B VSS:B EN:I IN0:B IN1:B OUT:B
x1 VDD ENB IN0 OUT VSS test_tg
x2 VDD EN IN1 OUT VSS test_tg
x3 VDD EN ENB VSS biasgen_inverter
.ends

* expanding   symbol:  libs/core_test/test_tg/test_tg.sym # of pins=5
** sym_path: /foss/designs/libs/core_test/test_tg/test_tg.sym
** sch_path: /foss/designs/libs/core_test/test_tg/test_tg.sch
.subckt test_tg VDD EN VIN VOUT VSS
*.PININFO VIN:B VOUT:B EN:I VDD:B VSS:B
XMTG1 VIN EN VOUT VSS nfet_05v0 L=0.60u W=1.5u nf=1 m=2
XMTG2 VOUT ENB VIN VDD pfet_05v0 L=0.50u W=1.5u nf=1 m=6
x1 VDD ENB EN VSS test_inv
.ends


* expanding   symbol:  libs/core_biasgen/biasgen_inverter/biasgen_inverter.sym # of pins=4
** sym_path: /foss/designs/libs/core_biasgen/biasgen_inverter/biasgen_inverter.sym
** sch_path: /foss/designs/libs/core_biasgen/biasgen_inverter/biasgen_inverter.sch
.subckt biasgen_inverter VDD IN OUT VSS
*.PININFO VDD:B VSS:B IN:I OUT:O
XMINV1 OUT IN VSS VSS nfet_05v0 L=0.60u W=0.42u nf=1 m=1
XMINV2 OUT IN VDD VDD pfet_05v0 L=0.50u W=0.60u nf=1 m=1
.ends


* expanding   symbol:  libs/core_test/test_inv/test_inv.sym # of pins=4
** sym_path: /foss/designs/libs/core_test/test_inv/test_inv.sym
** sch_path: /foss/designs/libs/core_test/test_inv/test_inv.sch
.subckt test_inv VDD OUT IN VSS
*.PININFO OUT:O IN:I VDD:B VSS:B
XMINV1 OUT IN VSS VSS nfet_05v0 L=0.60u W=0.42u nf=1 m=1
XMINV2 OUT IN VDD VDD pfet_05v0 L=0.50u W=0.60u nf=1 m=1
.ends

