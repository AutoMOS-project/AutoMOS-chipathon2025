* Extracted by KLayout with GF180 LVS runset on : 17/08/2025 21:25

.SUBCKT top_io PAD DVSS|VMINUS|VSS DVDD|VDD|VPLUS VSS DVDD DVSS
+ NDRIVE_X|ndrive_x_<1> NDRIVE_Y|ndrive_Y_<1> NDRIVE_X|ndrive_x_<2>
+ NDRIVE_Y|ndrive_y_<2> NDRIVE_X|ndrive_x_<3> NDRIVE_Y|ndrive_Y_<3>
+ NDRIVE_X|ndrive_x_<0> DVDD|VPLUS DVSS|VMINUS PDRIVE_X|pdrive_x_<0>
+ PDRIVE_Y|pdrive_y_<1> PDRIVE_X|pdrive_x_<1> PDRIVE_X|pdrive_x_<2>
+ PDRIVE_Y|pdrive_y_<2> PDRIVE_Y|pdrive_y_<3> PDRIVE_X|pdrive_x_<3>
+ NDRIVE_Y|ndrive_y_<0> PDRIVE_Y|pdrive_y_<0> SL|Z ENB EN A|AB SLB|ZB A|OE|PDRV
+ VRC PDRV|VDD A|IP_IN|PAD A|PDB_OUT|Z A|PUB_OUT|Z B|PD|PD_IN A|PU A|B|Z PU_B|Z
+ PD|ZB A|Z Y Z CS|Z IE|Z A|CS|IE ZB A|CS|OE|PDRV A|IE ASIG5V NDRIVE_X NDRIVE_Y
+ PDRIVE_X PDRIVE_Y PDRV|PDRV0 OE PDRV|PDRV1 A|SL A PDRV A|CS vss
M$1 DVDD \$114 NDRIVE_Y|ndrive_y_<0> DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$3 NDRIVE_X|ndrive_x_<0> SL|Z NDRIVE_Y|ndrive_y_<0> DVDD pfet_06v0 L=0.7U
+ W=72U AS=18.72P AD=25.2P PS=75.12U PD=112.2U
M$5 \$114 ENB \$113 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$6 DVDD EN \$114 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$7 \$114 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$8 PDRIVE_Y|pdrive_y_<0> \$113 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$10 PDRIVE_X|pdrive_x_<0> \$113 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$12 PDRIVE_X|pdrive_x_<1> \$120 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$14 PDRIVE_Y|pdrive_y_<1> \$120 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$16 DVDD A|AB \$119 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$17 \$119 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$18 \$120 ENB \$119 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$19 NDRIVE_X|ndrive_x_<1> SL|Z NDRIVE_Y|ndrive_Y_<1> DVDD pfet_06v0 L=0.7U
+ W=72U AS=25.2P AD=18.72P PS=112.2U PD=75.12U
M$21 DVDD \$119 NDRIVE_Y|ndrive_Y_<1> DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$23 DVDD \$125 NDRIVE_Y|ndrive_y_<2> DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$25 NDRIVE_X|ndrive_x_<2> SL|Z NDRIVE_Y|ndrive_y_<2> DVDD pfet_06v0 L=0.7U
+ W=72U AS=18.72P AD=25.2P PS=75.12U PD=112.2U
M$27 \$125 ENB \$124 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$28 DVDD EN \$125 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$29 \$125 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$30 PDRIVE_Y|pdrive_y_<2> \$124 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$32 PDRIVE_X|pdrive_x_<2> \$124 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$34 PDRIVE_X|pdrive_x_<3> \$130 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$36 PDRIVE_Y|pdrive_y_<3> \$130 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$38 DVDD A|AB \$129 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$39 \$129 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$40 \$130 ENB \$129 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$41 NDRIVE_X|ndrive_x_<3> SL|Z NDRIVE_Y|ndrive_Y_<3> DVDD pfet_06v0 L=0.7U
+ W=72U AS=25.2P AD=18.72P PS=112.2U PD=75.12U
M$43 DVDD \$129 NDRIVE_Y|ndrive_Y_<3> DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$45 DVDD \$138 NDRIVE_Y|ndrive_y_<0> DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$49 \$138 ENB \$137 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$50 DVDD EN \$138 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$51 \$138 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$52 PDRIVE_Y|pdrive_y_<0> \$137 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$54 PDRIVE_X|pdrive_x_<0> \$137 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$56 PDRIVE_X|pdrive_x_<1> \$144 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$58 PDRIVE_Y|pdrive_y_<1> \$144 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$60 DVDD A|AB \$143 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$61 \$143 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$62 \$144 ENB \$143 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$65 DVDD \$143 NDRIVE_Y|ndrive_Y_<1> DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$67 DVDD \$149 NDRIVE_Y|ndrive_y_<2> DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$71 \$149 ENB \$148 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$72 DVDD EN \$149 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$73 \$149 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$74 PDRIVE_Y|pdrive_y_<2> \$148 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$76 PDRIVE_X|pdrive_x_<2> \$148 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$78 PDRIVE_X|pdrive_x_<3> \$154 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$80 PDRIVE_Y|pdrive_y_<3> \$154 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$82 DVDD A|AB \$153 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$83 \$153 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$84 \$154 ENB \$153 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$87 DVDD \$153 NDRIVE_Y|ndrive_Y_<3> DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$89 \$241 VRC DVDD|VDD|VPLUS DVDD|VDD|VPLUS pfet_06v0 L=0.7U W=20U AS=6.1P
+ AD=5.2P PS=27.44U PD=22.08U
M$93 \$243 \$241 DVDD|VDD|VPLUS DVDD|VDD|VPLUS pfet_06v0 L=0.7U W=15U AS=3.9P
+ AD=4.8P PS=16.56U PD=21.92U
M$96 \$62 \$243 DVDD|VDD|VPLUS DVDD|VDD|VPLUS pfet_06v0 L=0.7U W=120U AS=32.1P
+ AD=32.1P PS=137.84U PD=137.84U
M$120 \$220 VRC DVDD|VPLUS DVDD|VPLUS pfet_06v0 L=0.7U W=20U AS=6.1P AD=5.2P
+ PS=27.44U PD=22.08U
M$124 \$222 \$220 DVDD|VPLUS DVDD|VPLUS pfet_06v0 L=0.7U W=15U AS=3.9P AD=4.8P
+ PS=16.56U PD=21.92U
M$127 \$59 \$222 DVDD|VPLUS DVDD|VPLUS pfet_06v0 L=0.7U W=120U AS=32.1P
+ AD=32.1P PS=137.84U PD=137.84U
M$151 NDRIVE_Y|ndrive_y_<0> DVSS NDRIVE_X|ndrive_x_<0> DVDD pfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$152 NDRIVE_X|ndrive_x_<1> DVSS NDRIVE_Y|ndrive_Y_<1> DVDD pfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$153 NDRIVE_Y|ndrive_y_<2> DVSS NDRIVE_X|ndrive_x_<2> DVDD pfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$154 NDRIVE_X|ndrive_x_<3> DVSS NDRIVE_Y|ndrive_Y_<3> DVDD pfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$155 \$258 A|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=2.1P
+ PS=10.4U PD=10.4U
M$158 DVDD \$258 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$159 ENB EN DVDD DVDD pfet_06v0 L=0.7U W=72U AS=23.04P AD=27.36P PS=103.68U
+ PD=129.12U
M$161 EN \$262 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$162 \$262 A|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=2.1P
+ PS=10.4U PD=10.4U
M$164 \$266 PDRV|VDD PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$165 PDRV|VDD A|OE|PDRV \$266 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$167 DVDD \$266 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$170 DVDD \$269 A|AB DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$171 \$269 \$271 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$172 \$271 A|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=2.1P
+ PS=10.4U PD=10.4U
M$174 \$274 A|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$175 SL|Z \$274 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$177 SLB|ZB SL|Z DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P PS=28.16U
+ PD=41.6U
M$180 \$323 A|CS|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=6U AS=2.1P
+ AD=2.1P PS=10.4U PD=10.4U
M$182 DVDD \$323 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$185 EN \$327 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$186 \$327 A|CS|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=6U AS=2.1P
+ AD=2.1P PS=10.4U PD=10.4U
M$188 \$331 PDRV|VDD PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$189 PDRV|VDD A|CS|OE|PDRV \$331 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P
+ AD=1.32P PS=3.52U PD=6.88U
M$190 DVDD \$331 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$192 DVDD \$334 A|AB DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$193 \$334 \$336 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$194 \$595 A|Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$195 \$336 A|CS|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=6U AS=2.1P
+ AD=2.1P PS=10.4U PD=10.4U
M$197 \$520 PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$198 \$341 A|CS|OE|PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$199 A|PDB_OUT|Z B|PD|PD_IN PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=12U AS=5.28P
+ AD=3.12P PS=27.52U PD=14.08U
M$200 PDRV|VDD A|B|Z A|PDB_OUT|Z PDRV|VDD pfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=5.28P PS=14.08U PD=27.52U
M$201 Y Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=84U AS=24.36P AD=24.36P
+ PS=111.92U PD=111.92U
M$207 \$522 B|PD|PD_IN PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$208 SL|Z \$341 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$212 A|B|Z \$522 \$517 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$213 A|PUB_OUT|Z A|B|Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=12U AS=5.28P
+ AD=3.12P PS=27.52U PD=14.08U
M$214 PDRV|VDD A|PU A|PUB_OUT|Z PDRV|VDD pfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=5.28P PS=14.08U PD=27.52U
M$215 A|PU B|PD|PD_IN A|B|Z PDRV|VDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=5.28P
+ PS=27.52U PD=27.52U
M$216 PDRV|VDD A|PU \$517 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$217 \$582 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U
+ PD=13.4U
M$219 \$576 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.05P AD=1.05P PS=5.9U
+ PD=5.9U
M$221 A|Z IE|Z DVDD DVDD pfet_06v0 L=0.7U W=24U AS=7.68P AD=7.68P PS=39.68U
+ PD=39.68U
M$224 DVDD A|IP_IN|PAD \$565 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P
+ PS=7.1U PD=7.1U
M$226 A|Z A|IP_IN|PAD \$565 DVDD pfet_06v0 L=0.7U W=4.3U AS=1.505P AD=1.505P
+ PS=7.85U PD=7.85U
M$228 DVSS \$576 \$565 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P PS=7.1U
+ PD=7.1U
M$230 A|Z \$582 \$576 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$231 \$578 \$582 A|Z DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$232 \$567 A|Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$233 \$497 PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$234 Z \$567 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=10U AS=3.05P AD=3.05P
+ PS=14.94U PD=14.94U
M$246 \$499 B|PD|PD_IN PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$247 A|B|Z \$499 \$495 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$251 PDRV|VDD A|PU \$495 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$252 \$634 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U
+ PD=13.4U
M$257 A|Z A|IP_IN|PAD \$593 DVDD pfet_06v0 L=0.7U W=4.3U AS=1.505P AD=1.505P
+ PS=7.85U PD=7.85U
M$259 \$612 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.05P AD=1.05P PS=5.9U
+ PD=5.9U
M$261 DVDD A|IP_IN|PAD \$593 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P
+ PS=7.1U PD=7.1U
M$263 DVSS \$612 \$593 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P PS=7.1U
+ PD=7.1U
M$265 A|Z \$634 \$612 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$266 \$614 \$634 A|Z DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$267 Z \$595 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=10U AS=3.05P AD=3.05P
+ PS=14.94U PD=14.94U
M$271 \$691 A|CS|IE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$272 PDRV|VDD A|CS|IE \$697 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$273 \$699 A|PDB_OUT|Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$274 PDRV|VDD A|PUB_OUT|Z \$705 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$275 IE|Z \$691 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$277 ZB IE|Z DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P PS=28.16U
+ PD=41.6U
M$279 ZB CS|Z DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P PS=41.6U
+ PD=28.16U
M$281 CS|Z \$697 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$283 Z \$699 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U PD=7.04U
M$285 PD|ZB Z DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P PS=28.16U
+ PD=41.6U
M$287 ZB PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P PS=41.6U
+ PD=28.16U
M$289 PU_B|Z \$705 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$291 \$744 A|IE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$292 IE|Z \$744 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$298 CS|Z \$750 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$300 PDRV|VDD A|CS|OE|PDRV \$750 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$301 \$752 A|PDB_OUT|Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$302 Z \$752 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U PD=7.04U
M$308 PU_B|Z \$758 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$310 PDRV|VDD A|PUB_OUT|Z \$758 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$311 DVDD \$1077 NDRIVE_Y|ndrive_y_<0> DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$315 \$1077 ENB \$1076 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$316 DVDD EN \$1077 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$317 \$1077 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$318 PDRIVE_Y|pdrive_y_<0> \$1076 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$320 PDRIVE_X|pdrive_x_<0> \$1076 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$322 PDRIVE_X|pdrive_x_<1> \$1083 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$324 PDRIVE_Y|pdrive_y_<1> \$1083 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$326 DVDD A|AB \$1082 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$327 \$1082 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$328 \$1083 ENB \$1082 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$331 DVDD \$1082 NDRIVE_Y|ndrive_Y_<1> DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$333 DVDD \$1088 NDRIVE_Y|ndrive_y_<2> DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$337 \$1088 ENB \$1087 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$338 DVDD EN \$1088 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$339 \$1088 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$340 PDRIVE_Y|pdrive_y_<2> \$1087 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$342 PDRIVE_X|pdrive_x_<2> \$1087 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$344 PDRIVE_X|pdrive_x_<3> \$1093 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P
+ AD=6.24P PS=37.4U PD=25.04U
M$346 PDRIVE_Y|pdrive_y_<3> \$1093 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$348 DVDD A|AB \$1092 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$349 \$1092 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$350 \$1093 ENB \$1092 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$353 DVDD \$1092 NDRIVE_Y|ndrive_Y_<3> DVDD pfet_06v0 L=0.7U W=24U AS=6.24P
+ AD=8.4P PS=25.04U PD=37.4U
M$355 DVDD \$1120 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P
+ PS=37.4U PD=25.04U
M$357 NDRIVE_X SL|Z NDRIVE_Y DVDD pfet_06v0 L=0.7U W=96U AS=29.28P AD=29.28P
+ PS=124.88U PD=124.88U
M$359 \$1120 ENB \$1119 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$360 DVDD EN \$1120 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$361 \$1120 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$362 PDRIVE_Y \$1119 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P
+ PS=37.4U PD=25.04U
M$364 PDRIVE_X \$1119 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P
+ PS=25.04U PD=37.4U
M$366 PDRIVE_X \$1126 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P
+ PS=37.4U PD=25.04U
M$368 PDRIVE_Y \$1126 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P
+ PS=25.04U PD=37.4U
M$370 DVDD A|AB \$1125 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$371 \$1125 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$372 \$1126 ENB \$1125 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$375 DVDD \$1125 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P
+ PS=25.04U PD=37.4U
M$377 DVDD \$1131 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P
+ PS=37.4U PD=25.04U
M$381 \$1131 ENB \$1130 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$382 DVDD EN \$1131 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$383 \$1131 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$384 PDRIVE_Y \$1130 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P
+ PS=37.4U PD=25.04U
M$386 PDRIVE_X \$1130 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P
+ PS=25.04U PD=37.4U
M$388 PDRIVE_X \$1136 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=8.4P AD=6.24P
+ PS=37.4U PD=25.04U
M$390 PDRIVE_Y \$1136 DVDD DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P
+ PS=25.04U PD=37.4U
M$392 DVDD A|AB \$1135 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$393 \$1135 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$394 \$1136 ENB \$1135 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$397 DVDD \$1135 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=24U AS=6.24P AD=8.4P
+ PS=25.04U PD=37.4U
M$399 \$1232 PDRV|PDRV0 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=0.78P PS=6.88U PD=3.52U
M$400 PDRV|VDD OE \$1232 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$402 DVDD \$1232 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$405 EN \$1236 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$406 \$1236 OE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$407 PDRV|VDD PDRV|PDRV1 \$1236 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P
+ AD=1.32P PS=3.52U PD=6.88U
M$408 \$1240 PDRV|VDD PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$409 PDRV|VDD OE \$1240 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$411 DVDD \$1240 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$414 DVDD \$1243 A|AB DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$415 \$1243 \$1245 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$416 \$1245 A PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$417 PDRV|VDD OE \$1245 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$418 \$1248 A|SL PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$419 SL|Z \$1248 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$424 NDRIVE_Y DVSS NDRIVE_X DVDD pfet_06v0 L=0.7U W=4.8U AS=2.112P AD=2.112P
+ PS=13.12U PD=13.12U
M$425 DVDD \$1307 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$428 EN \$1311 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$430 DVDD \$1315 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$433 DVDD \$1318 A|AB DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$434 \$1318 \$1320 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$435 \$1323 A|SL PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$436 SL|Z \$1323 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$441 \$1437 PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$446 \$1307 PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$447 PDRV|VDD OE \$1307 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$448 \$1311 OE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$449 PDRV|VDD PDRV \$1311 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$450 \$1315 PDRV|VDD PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$451 PDRV|VDD OE \$1315 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$452 \$1320 A PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$453 PDRV|VDD OE \$1320 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$454 \$1439 B|PD|PD_IN PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$455 A|B|Z \$1439 \$1435 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$457 PDRV|VDD A|PU \$1435 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$458 \$1476 PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$461 \$1482 B|PD|PD_IN PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$462 A|B|Z \$1482 \$1477 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$466 PDRV|VDD A|PU \$1477 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$467 \$1500 A|Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$474 \$1512 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U
+ PD=13.4U
M$476 \$1504 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.05P AD=1.05P PS=5.9U
+ PD=5.9U
M$481 DVDD A|IP_IN|PAD \$1491 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P
+ PS=7.1U PD=7.1U
M$483 A|Z A|IP_IN|PAD \$1491 DVDD pfet_06v0 L=0.7U W=4.3U AS=1.505P AD=1.505P
+ PS=7.85U PD=7.85U
M$485 DVSS \$1504 \$1491 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P PS=7.1U
+ PD=7.1U
M$487 A|Z \$1512 \$1504 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$488 \$1510 \$1512 A|Z DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$489 Z \$1500 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=10U AS=3.05P AD=3.05P
+ PS=14.94U PD=14.94U
M$493 \$1596 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U
+ PD=13.4U
M$495 \$1574 CS|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.05P AD=1.05P PS=5.9U
+ PD=5.9U
M$500 DVDD A|IP_IN|PAD \$1555 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P
+ PS=7.1U PD=7.1U
M$502 A|Z A|IP_IN|PAD \$1555 DVDD pfet_06v0 L=0.7U W=4.3U AS=1.505P AD=1.505P
+ PS=7.85U PD=7.85U
M$504 DVSS \$1574 \$1555 DVDD pfet_06v0 L=0.7U W=3.8U AS=1.33P AD=1.33P PS=7.1U
+ PD=7.1U
M$506 \$1557 A|Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$513 \$1581 A|IE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$514 IE|Z \$1581 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$520 CS|Z \$1587 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$522 PDRV|VDD A|CS \$1587 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$523 \$1589 A|PDB_OUT|Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$524 Z \$1589 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$530 PU_B|Z \$1595 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$532 PDRV|VDD A|PUB_OUT|Z \$1595 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$533 A|Z \$1596 \$1574 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$534 \$1577 \$1596 A|Z DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$535 Z \$1557 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=10U AS=3.05P AD=3.05P
+ PS=14.94U PD=14.94U
M$539 \$1658 A|IE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$540 IE|Z \$1658 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$546 CS|Z \$1664 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$548 PDRV|VDD A|CS \$1664 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$549 \$1666 A|PDB_OUT|Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$550 Z \$1666 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=2.1P AD=1.56P PS=10.4U
+ PD=7.04U
M$556 PU_B|Z \$1672 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.1P PS=7.04U
+ PD=10.4U
M$558 PDRV|VDD A|PUB_OUT|Z \$1672 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$559 DVSS|VMINUS \$62 DVDD|VDD|VPLUS vss nfet_06v0 L=0.7U W=4000U AS=1076P
+ AD=1076P PS=4243.04U PD=4243.04U
M$579 DVDD|VPLUS \$59 DVSS|VMINUS|VSS vss nfet_06v0 L=0.7U W=4000U AS=1076P
+ AD=1076P PS=4243.04U PD=4243.04U
M$719 PDRIVE_X|pdrive_x_<0> DVDD PDRIVE_Y|pdrive_y_<0> vss nfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$720 PDRIVE_Y|pdrive_y_<1> DVDD PDRIVE_X|pdrive_x_<1> vss nfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$721 PDRIVE_X|pdrive_x_<2> DVDD PDRIVE_Y|pdrive_y_<2> vss nfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$722 PDRIVE_Y|pdrive_y_<3> DVDD PDRIVE_X|pdrive_x_<3> vss nfet_06v0 L=0.7U
+ W=3.6U AS=1.584P AD=1.584P PS=9.84U PD=9.84U
M$723 NDRIVE_X|ndrive_x_<0> \$114 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$725 NDRIVE_Y|ndrive_y_<0> \$114 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$727 \$113 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$728 \$114 EN \$113 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$729 DVSS A|AB \$113 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$730 PDRIVE_Y|pdrive_y_<0> \$113 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$732 PDRIVE_Y|pdrive_y_<0> SLB|ZB PDRIVE_X|pdrive_x_<0> vss nfet_06v0 L=0.7U
+ W=36U AS=12.6P AD=12.6P PS=58.2U PD=58.2U
M$734 PDRIVE_Y|pdrive_y_<1> SLB|ZB PDRIVE_X|pdrive_x_<1> vss nfet_06v0 L=0.7U
+ W=36U AS=12.6P AD=12.6P PS=58.2U PD=58.2U
M$736 PDRIVE_Y|pdrive_y_<1> \$120 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$738 \$120 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$739 \$120 EN \$119 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$740 DVSS ENB \$120 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$741 NDRIVE_Y|ndrive_Y_<1> \$119 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$743 NDRIVE_X|ndrive_x_<1> \$119 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$745 NDRIVE_X|ndrive_x_<2> \$125 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$747 NDRIVE_Y|ndrive_y_<2> \$125 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$749 \$124 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$750 \$125 EN \$124 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$751 DVSS A|AB \$124 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$752 PDRIVE_Y|pdrive_y_<2> \$124 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$754 PDRIVE_Y|pdrive_y_<2> SLB|ZB PDRIVE_X|pdrive_x_<2> vss nfet_06v0 L=0.7U
+ W=36U AS=12.6P AD=12.6P PS=58.2U PD=58.2U
M$756 PDRIVE_Y|pdrive_y_<3> SLB|ZB PDRIVE_X|pdrive_x_<3> vss nfet_06v0 L=0.7U
+ W=36U AS=12.6P AD=12.6P PS=58.2U PD=58.2U
M$758 PDRIVE_Y|pdrive_y_<3> \$130 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$760 \$130 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$761 \$130 EN \$129 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$762 DVSS ENB \$130 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$763 NDRIVE_Y|ndrive_Y_<3> \$129 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$765 NDRIVE_X|ndrive_x_<3> \$129 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$767 NDRIVE_X|ndrive_x_<0> \$138 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$769 NDRIVE_Y|ndrive_y_<0> \$138 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$771 \$137 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$772 \$138 EN \$137 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$773 DVSS A|AB \$137 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$774 PDRIVE_Y|pdrive_y_<0> \$137 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$782 PDRIVE_Y|pdrive_y_<1> \$144 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$784 \$144 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$785 \$144 EN \$143 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$786 DVSS ENB \$144 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$787 NDRIVE_Y|ndrive_Y_<1> \$143 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$789 NDRIVE_X|ndrive_x_<1> \$143 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$791 NDRIVE_X|ndrive_x_<2> \$149 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$793 NDRIVE_Y|ndrive_y_<2> \$149 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$795 \$148 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$796 \$149 EN \$148 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$797 DVSS A|AB \$148 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$798 PDRIVE_Y|pdrive_y_<2> \$148 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$806 PDRIVE_Y|pdrive_y_<3> \$154 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$808 \$154 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$809 \$154 EN \$153 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$810 DVSS ENB \$154 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$811 NDRIVE_Y|ndrive_Y_<3> \$153 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$813 NDRIVE_X|ndrive_x_<3> \$153 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$815 \$241 VRC DVSS|VMINUS vss nfet_06v0 L=0.7U W=5U AS=2.2P AD=2.2P PS=10.88U
+ PD=10.88U
M$816 \$243 \$241 DVSS|VMINUS vss nfet_06v0 L=0.7U W=30U AS=8.7P AD=7.8P
+ PS=38.48U PD=33.12U
M$822 \$62 \$243 DVSS|VMINUS vss nfet_06v0 L=0.7U W=30U AS=7.8P AD=8.7P
+ PS=33.12U PD=38.48U
M$828 \$220 VRC DVSS|VMINUS|VSS vss nfet_06v0 L=0.7U W=5U AS=2.2P AD=2.2P
+ PS=10.88U PD=10.88U
M$829 \$222 \$220 DVSS|VMINUS|VSS vss nfet_06v0 L=0.7U W=30U AS=8.7P AD=7.8P
+ PS=38.48U PD=33.12U
M$835 \$59 \$222 DVSS|VMINUS|VSS vss nfet_06v0 L=0.7U W=30U AS=7.8P AD=8.7P
+ PS=33.12U PD=38.48U
M$841 \$322 A|CS|OE|PDRV VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$842 \$323 A|CS|OE|PDRV \$322 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$843 DVSS \$323 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$844 ENB EN DVSS vss nfet_06v0 L=0.7U W=36U AS=11.52P AD=13.68P PS=55.68U
+ PD=69.12U
M$846 EN \$327 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$847 \$328 A|CS|OE|PDRV \$327 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$848 VSS A|CS|OE|PDRV \$328 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$849 \$330 PDRV|VDD VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$850 \$331 A|CS|OE|PDRV \$330 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$851 DVSS \$331 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$853 DVSS \$334 A|AB vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$854 \$334 \$336 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$855 \$337 A|CS|OE|PDRV \$336 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$856 VSS A|CS|OE|PDRV \$337 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$857 \$341 A|CS|OE|PDRV VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$858 SL|Z \$341 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$860 SLB|ZB SL|Z DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P PS=16.16U
+ PD=23.6U
M$862 \$257 A|OE|PDRV VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$863 \$258 A|OE|PDRV \$257 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$864 DVSS \$258 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$867 EN \$262 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$868 \$263 A|OE|PDRV \$262 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$869 VSS A|OE|PDRV \$263 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$870 \$265 PDRV|VDD VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$871 \$266 A|OE|PDRV \$265 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$872 DVSS \$266 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$874 DVSS \$269 A|AB vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$875 \$269 \$271 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$876 \$272 A|OE|PDRV \$271 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$877 VSS A|OE|PDRV \$272 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$878 \$274 A|OE|PDRV VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$879 \$433 B|PD|PD_IN A|PDB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$880 VSS A|B|Z \$433 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$881 SL|Z \$274 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$885 \$436 A|B|Z A|PUB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$886 VSS A|PU \$436 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$887 \$455 B|PD|PD_IN A|PDB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$888 VSS A|B|Z \$455 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$889 \$458 A|B|Z A|PUB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$890 VSS A|PU \$458 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$891 \$522 B|PD|PD_IN VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$892 A|B|Z B|PD|PD_IN \$517 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$893 A|PU \$522 A|B|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$894 VSS A|PU \$517 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$895 \$497 PD|ZB DVSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$896 \$499 B|PD|PD_IN VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$897 A|B|Z B|PD|PD_IN \$495 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$898 A|PU \$499 A|B|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$899 VSS A|PU \$495 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$900 \$520 PD|ZB DVSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$901 DVSS \$582 \$578 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$902 \$610 IE|Z DVSS vss nfet_06v0 L=0.7U W=16U AS=4.736P AD=4.736P PS=22.16U
+ PD=22.16U
M$907 A|Z CS|Z \$576 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$908 \$578 CS|Z A|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$909 DVSS A|Z \$567 vss nfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U PD=13.4U
M$911 \$582 CS|Z DVSS vss nfet_06v0 L=0.7U W=4U AS=1.4P AD=1.4P PS=7.4U PD=7.4U
M$913 \$610 A|IP_IN|PAD \$617 vss nfet_06v0 L=0.7U W=10.6U AS=3.233P AD=3.233P
+ PS=15.69U PD=15.69U
M$917 A|Z A|IP_IN|PAD \$617 vss nfet_06v0 L=0.7U W=12U AS=3.66P AD=3.66P
+ PS=17.44U PD=17.44U
M$921 \$617 \$578 DVDD vss nfet_06v0 L=0.7U W=1.3U AS=0.572P AD=0.572P PS=3.48U
+ PD=3.48U
M$922 Z \$567 VSS vss nfet_06v0 L=0.7U W=2.5U AS=0.875P AD=0.875P PS=5.15U
+ PD=5.15U
M$924 Y Z VSS vss nfet_06v0 L=0.7U W=36U AS=10.44P AD=10.44P PS=55.92U PD=55.92U
M$930 \$634 CS|Z DVSS vss nfet_06v0 L=0.7U W=4U AS=1.4P AD=1.4P PS=7.4U PD=7.4U
M$932 DVSS \$634 \$614 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$933 \$662 IE|Z DVSS vss nfet_06v0 L=0.7U W=16U AS=4.736P AD=4.736P PS=22.16U
+ PD=22.16U
M$938 \$662 A|IP_IN|PAD \$664 vss nfet_06v0 L=0.7U W=10.6U AS=3.233P AD=3.233P
+ PS=15.69U PD=15.69U
M$942 A|Z A|IP_IN|PAD \$664 vss nfet_06v0 L=0.7U W=12U AS=3.66P AD=3.66P
+ PS=17.44U PD=17.44U
M$946 \$664 \$614 DVDD vss nfet_06v0 L=0.7U W=1.3U AS=0.572P AD=0.572P PS=3.48U
+ PD=3.48U
M$947 A|Z CS|Z \$612 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$948 \$614 CS|Z A|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$949 DVSS A|Z \$595 vss nfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U PD=13.4U
M$951 Z \$595 VSS vss nfet_06v0 L=0.7U W=2.5U AS=0.875P AD=0.875P PS=5.15U
+ PD=5.15U
M$959 \$744 A|IE VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$960 IE|Z \$744 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$962 ZB IE|Z DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P PS=16.16U
+ PD=23.6U
M$964 ZB CS|Z DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P AD=3.12P PS=23.6U
+ PD=16.16U
M$966 CS|Z \$750 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$968 VSS A|CS|OE|PDRV \$750 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$969 \$752 A|PDB_OUT|Z VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$970 Z \$752 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U PD=4.04U
M$972 PD|ZB Z DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P PS=16.16U
+ PD=23.6U
M$974 ZB PU_B|Z DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P AD=3.12P PS=23.6U
+ PD=16.16U
M$976 PU_B|Z \$758 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$978 VSS A|PUB_OUT|Z \$758 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$979 \$691 A|CS|IE VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$980 IE|Z \$691 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$986 CS|Z \$697 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$988 VSS A|CS|IE \$697 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$989 \$699 A|PDB_OUT|Z VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$990 Z \$699 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U PD=4.04U
M$996 PU_B|Z \$705 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$998 VSS A|PUB_OUT|Z \$705 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1003 NDRIVE_X|ndrive_x_<0> \$1077 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$1005 NDRIVE_Y|ndrive_y_<0> \$1077 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$1007 \$1076 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1008 \$1077 EN \$1076 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1009 DVSS A|AB \$1076 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1010 PDRIVE_Y|pdrive_y_<0> \$1076 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$1016 PDRIVE_Y|pdrive_y_<1> \$1083 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$1018 \$1083 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1019 \$1083 EN \$1082 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1020 DVSS ENB \$1083 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1021 NDRIVE_Y|ndrive_Y_<1> \$1082 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$1023 NDRIVE_X|ndrive_x_<1> \$1082 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$1025 NDRIVE_X|ndrive_x_<2> \$1088 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$1027 NDRIVE_Y|ndrive_y_<2> \$1088 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$1029 \$1087 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1030 \$1088 EN \$1087 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1031 DVSS A|AB \$1087 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1032 PDRIVE_Y|pdrive_y_<2> \$1087 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$1038 PDRIVE_Y|pdrive_y_<3> \$1093 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P
+ AD=3.12P PS=19.4U PD=13.04U
M$1040 \$1093 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1041 \$1093 EN \$1092 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1042 DVSS ENB \$1093 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1043 NDRIVE_Y|ndrive_Y_<3> \$1092 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=3.12P PS=13.04U PD=13.04U
M$1045 NDRIVE_X|ndrive_x_<3> \$1092 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P
+ AD=4.2P PS=13.04U PD=19.4U
M$1047 NDRIVE_X \$1120 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P AD=3.12P
+ PS=19.4U PD=13.04U
M$1049 NDRIVE_Y \$1120 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=13.04U PD=13.04U
M$1051 \$1119 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1052 \$1120 EN \$1119 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1053 DVSS A|AB \$1119 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1054 PDRIVE_Y \$1119 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P
+ PS=13.04U PD=19.4U
M$1056 PDRIVE_Y SLB|ZB PDRIVE_X vss nfet_06v0 L=0.7U W=48U AS=16.8P AD=16.8P
+ PS=77.6U PD=77.6U
M$1058 PDRIVE_X DVDD PDRIVE_Y vss nfet_06v0 L=0.7U W=4.8U AS=2.112P AD=2.112P
+ PS=13.12U PD=13.12U
M$1062 PDRIVE_Y \$1126 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P AD=3.12P
+ PS=19.4U PD=13.04U
M$1064 \$1126 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1065 \$1126 EN \$1125 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1066 DVSS ENB \$1126 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1067 NDRIVE_Y \$1125 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=13.04U PD=13.04U
M$1069 NDRIVE_X \$1125 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P
+ PS=13.04U PD=19.4U
M$1071 NDRIVE_X \$1131 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P AD=3.12P
+ PS=19.4U PD=13.04U
M$1073 NDRIVE_Y \$1131 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=13.04U PD=13.04U
M$1075 \$1130 ENB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1076 \$1131 EN \$1130 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1077 DVSS A|AB \$1130 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1078 PDRIVE_Y \$1130 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P
+ PS=13.04U PD=19.4U
M$1086 PDRIVE_Y \$1136 DVSS vss nfet_06v0 L=0.7U W=12U AS=4.2P AD=3.12P
+ PS=19.4U PD=13.04U
M$1088 \$1136 A|AB DVSS vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$1089 \$1136 EN \$1135 vss nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$1090 DVSS ENB \$1136 vss nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$1091 NDRIVE_Y \$1135 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=13.04U PD=13.04U
M$1093 NDRIVE_X \$1135 DVSS vss nfet_06v0 L=0.7U W=12U AS=3.12P AD=4.2P
+ PS=13.04U PD=19.4U
M$1095 \$1231 PDRV|PDRV0 VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$1096 \$1232 OE \$1231 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1097 DVSS \$1232 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1100 EN \$1236 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1101 \$1237 OE \$1236 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1102 VSS PDRV|PDRV1 \$1237 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$1103 \$1239 PDRV|VDD VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1104 \$1240 OE \$1239 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1105 DVSS \$1240 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1107 DVSS \$1243 A|AB vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1108 \$1243 \$1245 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1109 \$1246 A \$1245 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1110 VSS OE \$1246 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1111 \$1248 A|SL VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1112 SL|Z \$1248 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$1116 \$1306 PDRV VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1117 \$1307 OE \$1306 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1118 DVSS \$1307 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1121 EN \$1311 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1122 \$1312 OE \$1311 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1123 VSS PDRV \$1312 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1124 \$1314 PDRV|VDD VSS vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1125 \$1315 OE \$1314 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1126 DVSS \$1315 EN vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1128 DVSS \$1318 A|AB vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1129 \$1318 \$1320 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1130 \$1321 A \$1320 vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$1131 VSS OE \$1321 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1132 \$1323 A|SL VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1133 SL|Z \$1323 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$1137 \$1437 PD|ZB DVSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1138 \$1385 B|PD|PD_IN A|PDB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=0.78P PS=6.88U PD=3.52U
M$1139 VSS A|B|Z \$1385 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1140 \$1439 B|PD|PD_IN VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1141 A|B|Z B|PD|PD_IN \$1435 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1142 \$1388 A|B|Z A|PUB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$1143 VSS A|PU \$1388 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1144 A|PU \$1439 A|B|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1145 VSS A|PU \$1435 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1146 \$1430 B|PD|PD_IN A|PDB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=0.78P PS=6.88U PD=3.52U
M$1147 VSS A|B|Z \$1430 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1148 \$1482 B|PD|PD_IN VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1149 A|B|Z B|PD|PD_IN \$1477 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1150 \$1433 A|B|Z A|PUB_OUT|Z vss nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$1151 VSS A|PU \$1433 vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$1152 A|PU \$1482 A|B|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1153 VSS A|PU \$1477 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1154 A|Z CS|Z \$1504 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1155 \$1510 CS|Z A|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1156 DVSS A|Z \$1500 vss nfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U
+ PD=13.4U
M$1158 \$1476 PD|ZB DVSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1159 DVSS \$1512 \$1510 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1160 \$1528 IE|Z DVSS vss nfet_06v0 L=0.7U W=16U AS=4.736P AD=4.736P
+ PS=22.16U PD=22.16U
M$1165 \$1528 A|IP_IN|PAD \$1530 vss nfet_06v0 L=0.7U W=10.6U AS=3.233P
+ AD=3.233P PS=15.69U PD=15.69U
M$1169 A|Z A|IP_IN|PAD \$1530 vss nfet_06v0 L=0.7U W=12U AS=3.66P AD=3.66P
+ PS=17.44U PD=17.44U
M$1173 \$1530 \$1510 DVDD vss nfet_06v0 L=0.7U W=1.3U AS=0.572P AD=0.572P
+ PS=3.48U PD=3.48U
M$1174 \$1512 CS|Z DVSS vss nfet_06v0 L=0.7U W=4U AS=1.4P AD=1.4P PS=7.4U
+ PD=7.4U
M$1176 \$1581 A|IE VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1177 IE|Z \$1581 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$1183 CS|Z \$1587 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$1185 VSS A|CS \$1587 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1186 \$1589 A|PDB_OUT|Z VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1187 Z \$1589 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$1191 Z \$1500 VSS vss nfet_06v0 L=0.7U W=2.5U AS=0.875P AD=0.875P PS=5.15U
+ PD=5.15U
M$1195 PU_B|Z \$1595 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$1203 VSS A|PUB_OUT|Z \$1595 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1204 \$1596 CS|Z DVSS vss nfet_06v0 L=0.7U W=4U AS=1.4P AD=1.4P PS=7.4U
+ PD=7.4U
M$1206 DVSS \$1596 \$1577 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1207 \$1612 IE|Z DVSS vss nfet_06v0 L=0.7U W=16U AS=4.736P AD=4.736P
+ PS=22.16U PD=22.16U
M$1212 \$1612 A|IP_IN|PAD \$1616 vss nfet_06v0 L=0.7U W=10.6U AS=3.233P
+ AD=3.233P PS=15.69U PD=15.69U
M$1216 A|Z A|IP_IN|PAD \$1616 vss nfet_06v0 L=0.7U W=12U AS=3.66P AD=3.66P
+ PS=17.44U PD=17.44U
M$1220 \$1616 \$1577 DVDD vss nfet_06v0 L=0.7U W=1.3U AS=0.572P AD=0.572P
+ PS=3.48U PD=3.48U
M$1221 A|Z CS|Z \$1574 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1222 \$1577 CS|Z A|Z vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1223 DVSS A|Z \$1557 vss nfet_06v0 L=0.7U W=8U AS=2.8P AD=2.8P PS=13.4U
+ PD=13.4U
M$1225 \$1658 A|IE VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1226 IE|Z \$1658 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$1232 CS|Z \$1664 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$1234 VSS A|CS \$1664 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$1235 \$1666 A|PDB_OUT|Z VSS vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$1236 Z \$1666 DVSS vss nfet_06v0 L=0.7U W=3U AS=1.05P AD=0.78P PS=5.9U
+ PD=4.04U
M$1240 Z \$1557 VSS vss nfet_06v0 L=0.7U W=2.5U AS=0.875P AD=0.875P PS=5.15U
+ PD=5.15U
M$1244 PU_B|Z \$1672 DVSS vss nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.05P PS=4.04U
+ PD=5.9U
M$1252 VSS A|PUB_OUT|Z \$1672 vss nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
D$1253 VSS A|OE|PDRV diode_pd2nw_06v0 A=1.152P P=9.6U
D$1257 VSS PDRV|VDD diode_pd2nw_06v0 A=0.9216P P=7.68U
D$1259 VSS A|CS|OE|PDRV diode_pd2nw_06v0 A=1.152P P=9.6U
D$1265 A|OE|PDRV PDRV|VDD diode_pd2nw_06v0 A=2P P=8U
D$1267 A|CS|OE|PDRV PDRV|VDD diode_pd2nw_06v0 A=3P P=12U
D$1269 A|IP_IN|PAD DVDD diode_pd2nw_06v0 A=160P P=336U
D$1273 A|PU PDRV|VDD diode_pd2nw_06v0 A=4P P=16U
D$1274 B|PD|PD_IN PDRV|VDD diode_pd2nw_06v0 A=4P P=16U
D$1275 A|CS|IE PDRV|VDD diode_pd2nw_06v0 A=2P P=8U
D$1280 A|IE PDRV|VDD diode_pd2nw_06v0 A=3P P=12U
D$1281 ASIG5V DVDD diode_pd2nw_06v0 A=600P P=424U
D$1285 VSS PDRV|PDRV0 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$1286 VSS OE diode_pd2nw_06v0 A=1.3824P P=11.52U
D$1288 VSS PDRV|PDRV1 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$1291 VSS PDRV diode_pd2nw_06v0 A=0.4608P P=3.84U
D$1297 A PDRV|VDD diode_pd2nw_06v0 A=2P P=8U
D$1298 A|SL PDRV|VDD diode_pd2nw_06v0 A=2P P=8U
D$1307 A|CS PDRV|VDD diode_pd2nw_06v0 A=2P P=8U
R$1317 A|IP_IN|PAD \$520 vss 119393.75 ppolyf_u L=272.9U W=0.8U
R$1321 PAD A|IP_IN|PAD vss 24.5 ppolyf_u L=2.8U W=40U
R$1329 A|IP_IN|PAD \$497 vss 119393.75 ppolyf_u L=272.9U W=0.8U
R$1356 PDRV|VDD A|CS|IE vss 1706.25 ppolyf_u L=3.9U W=0.8U
R$1357 VSS A|OE|PDRV vss 1706.25 ppolyf_u L=3.9U W=0.8U
R$1361 DVDD|VPLUS VRC vss 335238.75 ppolyf_u L=766.26U W=0.8U
R$1362 DVDD|VDD|VPLUS VRC vss 335238.75 ppolyf_u L=766.26U W=0.8U
R$1363 PDRV|VDD A|IE vss 1706.25 ppolyf_u L=3.9U W=0.8U
R$1364 VSS A|CS|OE|PDRV vss 1706.25 ppolyf_u L=3.9U W=0.8U
R$1370 \$1437 A|IP_IN|PAD vss 119393.75 ppolyf_u L=272.9U W=0.8U
R$1381 A|IP_IN|PAD \$1476 vss 119393.75 ppolyf_u L=272.9U W=0.8U
R$1389 PDRV|VDD PDRV vss 350 ppolyf_u L=1.6U W=1.6U
C$1391 VRC DVSS|VMINUS|VSS 4.6e-12 cap_nmos_06v0 A=2000P P=560U
C$1395 VRC DVSS|VMINUS 4.6e-12 cap_nmos_06v0 A=2000P P=560U
C$1399 DVDD DVSS 1.95477e-11 cap_nmos_06v0 A=8499P P=2794U
C$1431 DVDD|VDD|VPLUS DVSS|VMINUS 2.07e-12 cap_nmos_06v0 A=900P P=240U
C$1435 DVDD|VPLUS DVSS|VMINUS|VSS 2.07e-12 cap_nmos_06v0 A=900P P=240U
M$1501 PAD PDRIVE_X|pdrive_x_<0> DVDD DVDD pfet_06v0_dss L=0.7U W=240U AS=468P
+ AD=446.4P PS=383.4U PD=262.32U
M$1503 PAD PDRIVE_Y|pdrive_y_<0> DVDD DVDD pfet_06v0_dss L=0.7U W=120U AS=73.2P
+ AD=373.2P PS=123.66U PD=138.66U
M$1504 DVDD PDRIVE_Y|pdrive_y_<1> PAD DVDD pfet_06v0_dss L=0.7U W=120U
+ AS=373.2P AD=73.2P PS=138.66U PD=123.66U
M$1505 PAD PDRIVE_X|pdrive_x_<1> DVDD DVDD pfet_06v0_dss L=0.7U W=240U
+ AS=446.4P AD=446.4P PS=262.32U PD=262.32U
M$1507 PAD PDRIVE_X|pdrive_x_<2> DVDD DVDD pfet_06v0_dss L=0.7U W=240U
+ AS=446.4P AD=446.4P PS=262.32U PD=262.32U
M$1509 PAD PDRIVE_Y|pdrive_y_<2> DVDD DVDD pfet_06v0_dss L=0.7U W=120U AS=73.2P
+ AD=373.2P PS=123.66U PD=138.66U
M$1510 DVDD PDRIVE_Y|pdrive_y_<3> PAD DVDD pfet_06v0_dss L=0.7U W=120U
+ AS=373.2P AD=73.2P PS=138.66U PD=123.66U
M$1511 PAD PDRIVE_X|pdrive_x_<3> DVDD DVDD pfet_06v0_dss L=0.7U W=240U
+ AS=446.4P AD=468P PS=262.32U PD=383.4U
M$1537 PAD PDRIVE_X DVDD DVDD pfet_06v0_dss L=0.7U W=480U AS=903.6P AD=903.6P
+ PS=570.12U PD=570.12U
M$1539 PAD PDRIVE_Y DVDD DVDD pfet_06v0_dss L=0.7U W=240U AS=446.4P AD=446.4P
+ PS=254.88U PD=254.88U
M$1549 PAD NDRIVE_X|ndrive_x_<0> DVSS vss nfet_06v0_dss L=1.15U W=114U
+ AS=90.06P AD=468.54P PS=232.74U PD=138.66U
M$1550 DVSS NDRIVE_Y|ndrive_y_<0> PAD vss nfet_06v0_dss L=1.15U W=114U
+ AS=468.54P AD=69.54P PS=138.66U PD=117.66U
M$1551 PAD NDRIVE_X|ndrive_x_<1> DVSS vss nfet_06v0_dss L=1.15U W=114U
+ AS=69.54P AD=468.54P PS=117.66U PD=138.66U
M$1552 DVSS NDRIVE_Y|ndrive_Y_<1> PAD vss nfet_06v0_dss L=1.15U W=114U
+ AS=468.54P AD=69.54P PS=138.66U PD=117.66U
M$1553 PAD NDRIVE_X|ndrive_x_<2> DVSS vss nfet_06v0_dss L=1.15U W=114U
+ AS=69.54P AD=468.54P PS=117.66U PD=138.66U
M$1554 DVSS NDRIVE_Y|ndrive_y_<2> PAD vss nfet_06v0_dss L=1.15U W=114U
+ AS=468.54P AD=69.54P PS=138.66U PD=117.66U
M$1555 PAD NDRIVE_X|ndrive_x_<3> DVSS vss nfet_06v0_dss L=1.15U W=114U
+ AS=69.54P AD=468.54P PS=117.66U PD=138.66U
M$1556 DVSS NDRIVE_Y|ndrive_Y_<3> PAD vss nfet_06v0_dss L=1.15U W=114U
+ AS=468.54P AD=90.06P PS=138.66U PD=232.74U
M$1573 PAD NDRIVE_X DVSS vss nfet_06v0_dss L=0.8U W=148U AS=96.94P AD=608.28P
+ PS=190.24U PD=180.88U
M$1574 DVSS NDRIVE_Y PAD vss nfet_06v0_dss L=0.8U W=148U AS=608.28P AD=96.94P
+ PS=180.88U PD=190.24U
.ENDS top_io
