** sch_path: /foss/designs/libs/tb_ldo/tb_ldo/tb_ldo/tb_ldo_dc/tb_ldo_dc.sch
**.subckt tb_ldo_dc
* noconn #net1
RL out GND 1.8k m=1
V1 VDD GND 2
V2 vref GND 0.9
I0 VDD net2 10u
CL net3 GND 0.1u m=1
Resr out net3 0.2 m=1
x1 VDD vref out net2 net1 GND ldo
IL out1 GND 1m
* noconn #net4
V3 vref1 GND 0.9
I1 VDD net5 10u
CL1 net6 GND 0.1u m=1
Resr1 out1 net6 0.2 m=1
x2 VDD vref1 out1 net5 net4 GND ldo
**** begin user architecture code



.control
save all

** Dropout voltage simulation
dc V1 0 5 0.01

** Measurements
meas dc Vdd_min FIND v(vdd) WHEN v(out)=1.8 RISE=1
let Vdropout=Vdd_min-1.8
print Vdropout

** Plots
setplot dc1
let vout=v(out)
let vin=v(vdd)
plot vout vin

write tb_ldo_dc1.raw

** Line regulation simulation
dc V1 2 5 0.001

** Measurements
meas dc Vout_max MAX v(out)
meas dc Vout_min MIN v(out)
let DeltaVdd=5-2
let DeltaVout=Vout_max-Vout_min
let Line_reg=DeltaVout/DeltaVdd
print Line_reg

** Plots
setplot dc2
let vout=v(out)
plot vout

write tb_ldo_dc2.raw

** Load regulation simulation
dc IL 0 2m 0.01m

** Measurements
meas dc Vout_max MAX v(out1)
meas dc Vout_min MIN v(out1)
let DeltaVout = Vout_max-Vout_min
let DeltaIload = 0-2m
let Load_reg = abs(DeltaVout/DeltaIload)
let Load_reg_por = (DeltaVout/1.8)*100
print Load_reg
print Load_reg_por

** Plots
setplot dc3
let vout=v(out1)
plot vout

write tb_ldo_dc3.raw

.endc
* ngspice commands



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
* .lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_statistical
* ngspice commands

**** end user architecture code
**.ends

* expanding   symbol:  libs/core_ldo/ldo/ldo/ldo.sym # of pins=6
** sym_path: /foss/designs/libs/core_ldo/ldo/ldo/ldo.sym
** sch_path: /foss/designs/libs/core_ldo/ldo/ldo/ldo.sch
.subckt ldo VDD VREF VOUT IBIAS SUB VSS
*.iopin VDD
*.iopin VSS
*.iopin VOUT
*.iopin SUB
*.iopin VREF
*.iopin IBIAS
XMpass VOUT Vota VDD VDD pfet_05v0 L=0.50u W=100.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=5
* noconn SUB
x1 VDD VREF Vfb Vota IBIAS VSS OTA
XR1[9] Vr_fb1[9] VOUT VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[8] Vr_fb1[8] Vr_fb1[9] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[7] Vr_fb1[7] Vr_fb1[8] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[6] Vr_fb1[6] Vr_fb1[7] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[5] Vr_fb1[5] Vr_fb1[6] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[4] Vr_fb1[4] Vr_fb1[5] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[3] Vr_fb1[3] Vr_fb1[4] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[2] Vr_fb1[2] Vr_fb1[3] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[1] Vr_fb1[1] Vr_fb1[2] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR1[0] Vfb Vr_fb1[1] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[9] Vr_fb2[9] Vfb VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[8] Vr_fb2[8] Vr_fb2[9] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[7] Vr_fb2[7] Vr_fb2[8] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[6] Vr_fb2[6] Vr_fb2[7] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[5] Vr_fb2[5] Vr_fb2[6] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[4] Vr_fb2[4] Vr_fb2[5] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[3] Vr_fb2[3] Vr_fb2[4] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[2] Vr_fb2[2] Vr_fb2[3] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[1] Vr_fb2[1] Vr_fb2[2] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XR2[0] VSS Vr_fb2[1] VDD ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRc[29] Vr_mc[29] Vmc VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[28] Vr_mc[28] Vr_mc[29] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[27] Vr_mc[27] Vr_mc[28] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[26] Vr_mc[26] Vr_mc[27] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[25] Vr_mc[25] Vr_mc[26] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[24] Vr_mc[24] Vr_mc[25] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[23] Vr_mc[23] Vr_mc[24] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[22] Vr_mc[22] Vr_mc[23] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[21] Vr_mc[21] Vr_mc[22] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[20] Vr_mc[20] Vr_mc[21] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[19] Vr_mc[19] Vr_mc[20] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[18] Vr_mc[18] Vr_mc[19] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[17] Vr_mc[17] Vr_mc[18] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[16] Vr_mc[16] Vr_mc[17] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[15] Vr_mc[15] Vr_mc[16] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[14] Vr_mc[14] Vr_mc[15] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[13] Vr_mc[13] Vr_mc[14] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[12] Vr_mc[12] Vr_mc[13] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[11] Vr_mc[11] Vr_mc[12] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[10] Vr_mc[10] Vr_mc[11] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[9] Vr_mc[9] Vr_mc[10] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[8] Vr_mc[8] Vr_mc[9] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[7] Vr_mc[7] Vr_mc[8] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[6] Vr_mc[6] Vr_mc[7] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[5] Vr_mc[5] Vr_mc[6] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[4] Vr_mc[4] Vr_mc[5] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[3] Vr_mc[3] Vr_mc[4] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[2] Vr_mc[2] Vr_mc[3] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[1] Vr_mc[1] Vr_mc[2] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XRc[0] VOUT Vr_mc[1] VDD ppolyf_u_1k r_width=1e-6 r_length=10e-6 m=1
XCc Vota Vmc cap_mim_1f0fF c_width=25e-6 c_length=25e-6 m=4
XRfb_dummy_L[7] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[6] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[5] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[4] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[3] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[2] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[1] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_L[0] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[13] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[12] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[11] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[10] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[9] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[8] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[7] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[6] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[5] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[4] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[3] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[2] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[1] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
XRfb_dummy_TB[0] VSS VSS VSS ppolyf_u_1k r_width=1e-6 r_length=5e-6 m=1
.ends


* expanding   symbol:  libs/core_ldo/ldo/ldo_OTA/OTA.sym # of pins=6
** sym_path: /foss/designs/libs/core_ldo/ldo/ldo_OTA/OTA.sym
** sch_path: /foss/designs/libs/core_ldo/ldo/ldo_OTA/OTA.sch
.subckt OTA VDD VREF VFB VOTA IBIAS VSS
*.iopin VDD
*.iopin VSS
*.iopin VOTA
*.iopin VREF
*.iopin IBIAS
*.iopin VFB
XM3 net2 net2 VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net3 net3 VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net4 net2 VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 VOTA net3 VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=3
XM9 IBIAS IBIAS VSS VSS nfet_05v0 L=1.00u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM10 net1 IBIAS VSS VSS nfet_05v0 L=1.00u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net4 net4 VSS VSS nfet_05v0 L=1.00u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 VOTA net4 VSS VSS nfet_05v0 L=1.00u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=3
XM1 net2 VREF net1 VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 net3 VFB net1 VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_L[3] VDD VDD VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_L[2] VDD VDD VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_L[1] VDD VDD VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_L[0] VDD VDD VDD VDD pfet_05v0 L=1.00u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[9] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[8] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[7] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[6] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[5] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[4] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[3] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[2] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[1] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMpota_dummy_TB[0] VDD VDD VDD VDD pfet_05v0 L=0.50u W=11.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_L[1] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_L[0] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[7] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[6] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[5] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[4] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[3] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[2] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[1] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMndiff_dummy_TB[0] VSS VSS VSS VSS nfet_05v0 L=0.60u W=70.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_L[3] VSS VSS VSS VSS nfet_05v0 L=1.00u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_L[2] VSS VSS VSS VSS nfet_05v0 L=1.00u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_L[1] VSS VSS VSS VSS nfet_05v0 L=1.00u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_L[0] VSS VSS VSS VSS nfet_05v0 L=1.00u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[7] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[6] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[5] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[4] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[3] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[2] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[1] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnota_dummy_TB[0] VSS VSS VSS VSS nfet_05v0 L=0.60u W=2.50u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_L[1] VSS VSS VSS VSS nfet_05v0 L=1.00u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_L[0] VSS VSS VSS VSS nfet_05v0 L=1.00u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[7] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[6] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[5] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[4] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[3] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[2] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[1] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XMnbias_dummy_TB[0] VSS VSS VSS VSS nfet_05v0 L=0.60u W=6.00u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
