* NGSPICE file created from top_amux_2x1.ext - technology: gf180mcuD

.subckt top_amux_2x1 VDD VSS EN IN0 IN1 OUT
X0 IN1 a_n28035_n33468# OUT VDD pfet_05v0 ad=1.155p pd=4.54u as=1.155p ps=4.54u w=1.5u l=0.5u M=6
X1 OUT a_n28035_n31800# IN0 VSS nfet_05v0 ad=1.095p pd=4.46u as=1.095p ps=4.46u w=1.5u l=0.6u M=2
X2 IN0 a_n28035_n32634# OUT VDD pfet_05v0 ad=1.155p pd=4.54u as=1.155p ps=4.54u w=1.5u l=0.5u M=6
X3 OUT EN IN1 VSS nfet_05v0 ad=1.095p pd=4.46u as=1.095p ps=4.46u w=1.5u l=0.6u M=2
X4 VDD EN a_n28035_n33468# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X5 VDD EN a_n28035_n31800# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X6 VSS EN a_n28035_n31800# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X7 VDD a_n28035_n31800# a_n28035_n32634# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X8 VSS a_n28035_n31800# a_n28035_n32634# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X9 VSS EN a_n28035_n33468# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
.ends

