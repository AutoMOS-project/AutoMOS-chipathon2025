* NGSPICE file created from bandgap.ext - technology: gf180mcuD

.subckt cap_mim$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=16u c_length=16u
.ends

.subckt bandgap_opamp$1 VSS vn vp ibias VDD vout
Xcap_mim$1_0 a_n5609_n2907# vout cap_mim$1
X0 vout ibias VDD VDD pfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=1u M=8
X1 VDD VDD VDD VDD pfet_05v0 ad=1.16p pd=5.16u as=14.04p ps=76.32u w=2u l=1u M=4
X2 VSS VSS VSS VSS nfet_05v0 ad=0.29p pd=2.16u as=11.8p ps=87.2u w=0.5u l=2u M=10
X3 a_n3877_n280# ibias VDD VDD pfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=1u M=2
X4 vout a_n5609_n2907# VSS VSS nfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=2u M=16
X5 VDD VDD VDD VDD pfet_05v0 ad=0.29p pd=2.16u as=0 ps=0 w=0.5u l=1u M=2
X6 a_n5609_n2907# vp a_n3877_n280# VDD pfet_05v0 ad=1.2p pd=5.2u as=1.2p ps=5.2u w=2u l=1u M=2
X7 a_n6009_n3115# vn a_n3877_n280# VDD pfet_05v0 ad=1.2p pd=5.2u as=1.2p ps=5.2u w=2u l=1u M=2
X8 ibias ibias VDD VDD pfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=1u M=2
X9 a_n5609_n2907# a_n6009_n3115# VSS VSS nfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=2u M=2
X10 a_n6009_n3115# a_n6009_n3115# VSS VSS nfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=2u M=2
.ends

.subckt ppolyf_u_high_Rs_resistor$1 a_n128_0# a_1800_0# a_n352_0#
X0 a_n128_0# a_1800_0# a_n352_0# ppolyf_u_1k_6p0 r_width=1u r_length=9u
.ends

.subckt ppolyf_u_high_Rs_resistor a_900_0# a_n128_0# a_n352_0#
X0 a_n128_0# a_900_0# a_n352_0# ppolyf_u_1k_6p0 r_width=1u r_length=4.5u
.ends

.subckt bandgap vpref vpref_fb VSS VDD ICTAT VZTC IZTC VBG IPTAT
Xbandgap_opamp$1_0 VSS bandgap_opamp$1_0/vn bandgap_opamp$1_0/vp bandgap_opamp$1_0/ibias
+ VDD vpref_fb bandgap_opamp$1
Xppolyf_u_high_Rs_resistor$1_0[0|0] a_n22908_n917# m2_n28372_9003# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[1|0] m1_n25775_7400# m2_n28372_8203# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[2|0] m1_n25775_7400# m2_n28372_7403# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[3|0] m1_n25775_5800# m2_n28372_6603# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[4|0] m1_n25775_5800# m2_n28372_5803# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[5|0] m1_n25775_4200# m2_n28372_5003# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[6|0] m1_n25775_4200# m2_n28372_4203# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[7|0] m1_n25775_2600# m2_n28372_3403# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[8|0] m1_n25775_2600# m2_n28372_2603# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[9|0] m1_n25775_1000# m2_n28372_1803# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[10|0] m1_n25775_1000# m2_n28372_1003# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[11|0] VSS m2_n28372_203# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[0|1] m2_n28372_9003# m2_n30972_9003# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[1|1] m2_n28372_8203# m2_n30972_8203# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[2|1] m2_n28372_7403# m2_n30972_7403# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[3|1] m2_n28372_6603# m2_n30972_6603# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[4|1] m2_n28372_5803# m2_n30972_5803# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[5|1] m2_n28372_5003# m2_n30972_5003# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[6|1] m2_n28372_4203# m2_n30972_4203# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[7|1] m2_n28372_3403# m2_n30972_3403# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[8|1] m2_n28372_2603# m2_n30972_2603# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[9|1] m2_n28372_1803# m2_n30972_1803# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[10|1] m2_n28372_1003# m2_n30972_1003# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[11|1] m2_n28372_203# m2_n30972_203# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[0|2] m2_n30972_9003# m1_n32960_8202# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[1|2] m2_n30972_8203# m1_n32960_8202# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[2|2] m2_n30972_7403# m1_n32960_6602# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[3|2] m2_n30972_6603# m1_n32960_6602# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[4|2] m2_n30972_5803# m1_n32960_5002# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[5|2] m2_n30972_5003# m1_n32960_5002# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[6|2] m2_n30972_4203# m1_n32960_3402# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[7|2] m2_n30972_3403# m1_n32960_3402# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[8|2] m2_n30972_2603# m1_n32960_1802# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[9|2] m2_n30972_1803# m1_n32960_1802# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[10|2] m2_n30972_1003# m1_n32960_202# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor$1_0[11|2] m2_n30972_203# m1_n32960_202# VSS ppolyf_u_high_Rs_resistor$1
Xppolyf_u_high_Rs_resistor_0[0|0] m2_2232_15505# m1_1154_15445# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[1|0] m2_2232_16305# m1_1154_15445# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[0|1] m2_3831_15502# m2_2232_15505# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[1|1] m2_3831_16305# m2_2232_16305# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[0|2] m2_5433_15504# m2_3831_15502# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[1|2] m2_5432_16305# m2_3831_16305# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[0|3] m3_9250_15170# m2_5433_15504# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_0[1|3] m3_9499_6017# m2_5432_16305# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|0] m2_n6118_n11554# VSS VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|0] m2_n6118_n10554# m1_n7199_n10552# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|0] m2_n6118_n9554# m1_n7199_n10552# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|0] m2_n6118_n8554# m2_n9000_n8552# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|0] m2_n6118_n7554# VSS VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|1] m2_n4518_n11554# m2_n6118_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|1] m2_n4518_n10554# m2_n6118_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|1] m2_n4518_n9554# m2_n6118_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|1] m2_n4518_n8554# m2_n6118_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|1] m2_n4518_n7554# m2_n6118_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|2] m2_n2918_n11554# m2_n4518_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|2] m2_n2918_n10554# m2_n4518_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|2] m2_n2918_n9554# m2_n4518_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|2] m2_n2918_n8554# m2_n4518_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|2] m2_n2918_n7554# m2_n4518_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|3] m2_n1318_n11554# m2_n2918_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|3] m2_n1318_n10554# m2_n2918_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|3] m2_n1318_n9554# m2_n2918_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|3] m2_n1318_n8554# m2_n2918_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|3] m2_n1318_n7554# m2_n2918_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|4] m2_282_n11554# m2_n1318_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|4] m2_282_n10554# m2_n1318_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|4] m2_282_n9554# m2_n1318_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|4] m2_282_n8554# m2_n1318_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|4] m2_282_n7554# m2_n1318_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|5] m2_1882_n11554# m2_282_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|5] m2_1882_n10554# m2_282_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|5] m2_1882_n9554# m2_282_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|5] m2_1882_n8554# m2_282_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|5] m2_1882_n7554# m2_282_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|6] m2_3482_n11554# m2_1882_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|6] m2_3482_n10554# m2_1882_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|6] m2_3477_n9001# m2_1882_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|6] m2_3482_n8554# m2_1882_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|6] m2_3482_n7554# m2_1882_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|7] m2_5082_n11554# m2_3482_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|7] m2_5082_n10554# m2_3482_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|7] m2_5082_n9554# m1_4002_n9557# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|7] m2_5082_n8554# m2_3482_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|7] m2_5082_n7554# m2_3482_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|8] m2_6682_n11554# m2_5082_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|8] m2_6682_n10554# m2_5082_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|8] m2_6682_n9554# m2_5082_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|8] m2_6682_n8554# m2_5082_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|8] m2_6682_n7554# m2_5082_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|9] m2_8282_n11554# m2_6682_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|9] m2_8282_n10229# m2_6682_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|9] m2_8280_n9231# m2_6682_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|9] m2_8282_n8227# m2_6682_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|9] m2_8282_n7554# m2_6682_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|10] m2_9882_n11554# m2_8282_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|10] m2_9882_n10554# m2_8801_n9876# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|10] m2_9882_n9554# m1_8799_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|10] m2_9882_n8554# m1_8799_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|10] m2_9882_n7554# m2_8282_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|11] m2_11481_n11379# m2_9882_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|11] m2_12002_n11555# m2_9882_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|11] m2_11482_n9554# m2_9882_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|11] m2_11482_n8554# m2_9882_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|11] m2_11481_n7731# m2_9882_n7554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|12] m2_13082_n11554# m2_12002_n11555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|12] m2_13082_n10554# m2_11481_n11379# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|12] m2_13082_n9731# m2_11482_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|12] m2_11999_n7880# m2_11482_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|12] m2_13081_n7555# m2_11999_n7880# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|13] m2_14682_n11554# m2_13082_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|13] m2_14682_n10554# m2_13082_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|13] m2_14682_n9554# m2_8801_n9876# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|13] m2_14682_n8554# m2_11481_n7731# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|13] m2_14681_n7555# m2_13081_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|14] m2_16282_n11554# m2_14682_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|14] m2_13082_n9731# m2_14682_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|14] m1_16283_n9553# m2_14682_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|14] m1_16283_n9553# m2_14682_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|14] m2_16281_n7555# m2_14681_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|15] m2_17882_n11554# m2_16282_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|15] m2_17882_n10554# m2_8282_n10229# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|15] m2_17882_n9554# m2_8280_n9231# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|15] m2_17882_n8554# m2_8282_n8227# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|15] m2_17881_n7555# m2_16281_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|16] m2_19482_n11554# m2_17882_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|16] m2_19482_n10554# m2_17882_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|16] m2_19482_n9554# m2_17882_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|16] m2_19482_n8554# m2_17882_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|16] m2_19481_n7555# m2_17881_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|17] m2_21082_n11554# m2_19482_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|17] m2_21082_n10554# m2_19482_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|17] bandgap_opamp$1_0/vp m2_19482_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|17] m2_21082_n8554# m2_19482_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|17] m2_21081_n7555# m2_19481_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|18] m2_22682_n11554# m2_21082_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|18] m2_22682_n10554# m2_21082_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|18] m2_22682_n9554# m2_3477_n9001# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|18] m2_22682_n8554# m2_21082_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|18] m2_22681_n7555# m2_21081_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|19] m2_24282_n11554# m2_22682_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|19] m2_24282_n10554# m2_22682_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|19] m2_24282_n9554# m2_22682_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|19] m2_24282_n8554# m2_22682_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|19] m2_24281_n7555# m2_22681_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|20] m2_25882_n11554# m2_24282_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|20] m2_25882_n10554# m2_24282_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|20] m2_25882_n9554# m2_24282_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|20] m2_25882_n8554# m2_24282_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|20] m2_25881_n7555# m2_24281_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|21] m2_27482_n11554# m2_25882_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|21] m2_27482_n10554# m2_25882_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|21] m2_27482_n9554# m2_25882_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|21] m2_27482_n8554# m2_25882_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|21] m2_27481_n7555# m2_25881_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|22] m2_29082_n11554# m2_27482_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|22] m2_29082_n10554# m2_27482_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|22] m2_29082_n9554# m2_27482_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|22] m2_29082_n8554# m2_27482_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|22] m2_29081_n7555# m2_27481_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|23] m2_30682_n11554# m2_29082_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|23] m2_30682_n10554# m2_29082_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|23] m2_30682_n9554# m2_29082_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|23] m2_30682_n8554# m2_29082_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|23] m2_30681_n7555# m2_29081_n7555# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[0|24] VZTC m2_30682_n11554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[1|24] VBG m2_30682_n10554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[2|24] m1_32282_n9554# m2_30682_n9554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[3|24] m1_32282_n9554# m2_30682_n8554# VSS ppolyf_u_high_Rs_resistor
Xppolyf_u_high_Rs_resistor_1[4|24] w_11108_n5057# m2_30681_n7555# VSS ppolyf_u_high_Rs_resistor
X0 VSS VSS m1_4002_n9557# pnp_05p00x00p42 M=16
X1 a_n5453_5070# a_n7625_4860# a_n5733_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X2 a_n5453_5070# a_12938_n3515# a_12818_n3307# w_11108_n5057# nfet_05v0 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=0.6u M=16
X3 IZTC m3_9499_6017# a_11246_6327# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=6
X4 a_n22908_n917# a_n7625_4860# VDD VDD pfet_05v0 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=0.5u M=16
X5 a_n4727_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X6 VSS a_n22908_n917# VSS VSS nfet_05v0 ad=2.4p pd=9.2u as=0.10291n ps=0.43224m w=4u l=1u M=32
X7 IZTC a_n7625_4860# a_n7745_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X8 VSS a_n5453_5070# VSS VSS nfet_05v0 ad=2.4p pd=9.2u as=0 ps=0 w=4u l=1u M=32
X9 a_14264_6327# m3_9250_15170# VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=4
X10 VDD VDD VDD VDD pfet_05v0 ad=1.856p pd=7.56u as=0.25402n ps=0.97778m w=3.2u l=0.8u M=2
X11 VSS VSS VSS VSS nfet_05v0 ad=0.29p pd=2.16u as=0 ps=0 w=0.5u l=2u M=2
X12 VZTC m3_9499_6017# a_13258_6327# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=6
X13 VSS a_n22908_n917# a_n7625_4860# a_n7625_4860# pfet_05v0 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=0.5u M=32
X14 IPTAT a_n7625_4860# a_n3721_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X15 a_12938_n3515# a_12938_n3515# w_11108_n5057# w_11108_n5057# nfet_05v0 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=0.6u M=16
X16 VSS VSS a_12818_n3307# pnp_05p00x00p42 M=2
X17 VSS VSS VSS pnp_05p00x00p42 M=10
X18 a_n7745_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X19 a_n1669_n50# a_n3315_n258# VSS VSS nfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=2u M=2
X20 VSS a_n22908_n917# vpref vpref pfet_05v0 ad=2.4p pd=9.2u as=2.4p ps=9.2u w=4u l=0.5u M=32
X21 ICTAT m3_9499_6017# a_14264_6327# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=4
X22 m3_9250_15170# m3_9499_6017# a_16276_6327# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=4
X23 a_15270_6327# m3_9250_15170# VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=4
X24 VDD VDD VDD VDD pfet_05v0 ad=7.424p pd=26.76u as=0 ps=0 w=12.8u l=3.2u M=2
X25 VDD VDD VDD VDD pfet_05v0 ad=7.424p pd=26.76u as=0 ps=0 w=12.8u l=0.8u M=4
X26 a_n6739_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X27 VDD VDD VDD VDD pfet_05v0 ad=1.856p pd=7.56u as=0 ps=0 w=3.2u l=0.8u M=4
X28 a_n7625_4860# a_n3315_n258# VSS VSS nfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=2u M=2
X29 w_11108_n5057# w_11108_n5057# w_11108_n5057# w_11108_n5057# nfet_05v0 ad=2.32p pd=9.16u as=21.91862p ps=88.935u w=4u l=0.6u M=8
X30 a_n3315_n258# a_n3315_n258# VSS VSS nfet_05v0 ad=0.3p pd=2.2u as=0.3p ps=2.2u w=0.5u l=2u M=2
X31 a_16276_6327# m3_9250_15170# VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=4
X32 VSS VSS bandgap_opamp$1_0/vn pnp_05p00x00p42 M=2
X33 a_n703_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X34 VBG a_n7625_4860# a_n4727_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X35 VDD VDD VDD VDD pfet_05v0 ad=7.424p pd=26.76u as=0 ps=0 w=12.8u l=0.8u M=2
X36 a_12938_n3515# m3_9499_6017# a_15270_6327# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=4
X37 a_13258_6327# m3_9250_15170# VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=6
X38 VZTC a_n7625_4860# a_n6739_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X39 VSS VSS m2_n9000_n8552# pnp_05p00x00p42 M=2
X40 a_n3315_n258# a_n7625_4860# a_n2715_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X41 a_11246_6327# m3_9250_15170# VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=6
X42 a_n7625_4860# a_n7625_4860# VDD VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=3.2u M=2
X43 a_n1669_n50# a_n22908_n917# bandgap_opamp$1_0/ibias VSS nfet_05v0 ad=0.73p pd=3.46u as=0.73p ps=3.46u w=1u l=0.6u
X44 a_n2715_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X45 a_n3721_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X46 a_n1709_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X47 a_n5733_5070# vpref VDD VDD pfet_05v0 ad=1.92p pd=7.6u as=1.92p ps=7.6u w=3.2u l=0.8u M=2
X48 bandgap_opamp$1_0/vn a_n7625_4860# a_n703_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X49 bandgap_opamp$1_0/vp a_n7625_4860# a_n1709_5070# VDD pfet_05v0 ad=7.68p pd=26.8u as=7.68p ps=26.8u w=12.8u l=0.8u M=2
X50 VSS a_n5453_5070# m3_9499_6017# VSS nfet_05v0 ad=0.73p pd=3.46u as=0.73p ps=3.46u w=1u l=4u
.ends

