* Extracted by KLayout with GF180MCU LVS runset on : 01/09/2025 05:06

.SUBCKT bandgap I1_default_C I1_default_B I1_default_E SUB
M$1 \$858 \$945 \$857 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$2 \$860 \$946 \$859 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$3 \$862 \$947 \$861 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$4 \$864 \$948 \$863 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$5 \$866 \$949 \$865 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$6 \$868 \$950 \$867 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$7 \$870 \$951 \$869 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$8 \$872 \$952 \$871 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$9 \$842 \$937 \$841 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P PS=9.54U
+ PD=9.54U
M$10 \$844 \$938 \$843 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$11 \$846 \$939 \$845 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$12 \$848 \$940 \$847 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$13 \$850 \$941 \$849 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$14 \$852 \$942 \$851 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$15 \$854 \$943 \$853 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$16 \$856 \$944 \$855 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$17 \$962 \$1049 \$961 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$18 \$964 \$1050 \$963 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$19 \$966 \$1051 \$965 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$20 \$968 \$1052 \$967 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$21 \$970 \$1053 \$969 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$22 \$972 \$1054 \$971 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$23 \$974 \$1055 \$973 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$24 \$976 \$1056 \$975 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$25 \$978 \$993 \$977 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$26 \$980 \$994 \$979 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$27 \$982 \$995 \$981 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$28 \$984 \$996 \$983 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$29 \$986 \$997 \$985 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$30 \$988 \$998 \$987 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$31 \$990 \$999 \$989 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$32 \$992 \$1000 \$991 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$33 \$1082 \$1113 \$1081 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$34 \$1084 \$1114 \$1083 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$35 \$1086 \$1115 \$1085 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$36 \$1088 \$1116 \$1087 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$37 \$1090 \$1117 \$1089 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$38 \$1092 \$1118 \$1091 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$39 \$1094 \$1119 \$1093 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$40 \$1096 \$1120 \$1095 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$41 \$1098 \$1121 \$1097 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$42 \$1100 \$1122 \$1099 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$43 \$1102 \$1123 \$1101 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$44 \$1104 \$1124 \$1103 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$45 \$1106 \$1125 \$1105 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$46 \$1108 \$1126 \$1107 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$47 \$1110 \$1127 \$1109 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$48 \$1112 \$1128 \$1111 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$49 \$1162 \$1224 \$1161 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$50 \$1164 \$1225 \$1163 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$51 \$1166 \$1226 \$1165 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$52 \$1168 \$1227 \$1167 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$53 \$1170 \$1228 \$1169 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$54 \$1172 \$1229 \$1171 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$55 \$1174 \$1230 \$1173 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$56 \$1176 \$1231 \$1175 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$57 \$1178 \$1232 \$1177 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$58 \$1180 \$1233 \$1179 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$59 \$1182 \$1234 \$1181 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$60 \$1184 \$1235 \$1183 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$61 \$1186 \$1236 \$1185 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$62 \$1188 \$1237 \$1187 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$63 \$1190 \$1238 \$1189 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$64 \$1192 \$1239 \$1191 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$65 \$1267 \$1313 \$1266 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$66 \$1269 \$1314 \$1268 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$67 \$1271 \$1315 \$1270 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$68 \$1273 \$1316 \$1272 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$69 \$1275 \$1317 \$1274 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$70 \$1277 \$1318 \$1276 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$71 \$1279 \$1319 \$1278 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$72 \$1281 \$1320 \$1280 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$73 \$1283 \$1321 \$1282 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$74 \$1285 \$1322 \$1284 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$75 \$1287 \$1323 \$1286 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$76 \$1289 \$1324 \$1288 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$77 \$1291 \$1325 \$1290 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$78 \$1293 \$1326 \$1292 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$79 \$1295 \$1327 \$1294 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$80 \$1297 \$1328 \$1296 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$81 \$1402 \$1448 \$1401 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$82 \$1404 \$1449 \$1403 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$83 \$1406 \$1450 \$1405 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$84 \$1408 \$1451 \$1407 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$85 \$1410 \$1452 \$1409 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$86 \$1412 \$1453 \$1411 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$87 \$1414 \$1454 \$1413 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$88 \$1416 \$1455 \$1415 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$89 \$1418 \$1456 \$1417 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$90 \$1420 \$1457 \$1419 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$91 \$1422 \$1458 \$1421 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$92 \$1424 \$1459 \$1423 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$93 \$1426 \$1460 \$1425 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$94 \$1428 \$1461 \$1427 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$95 \$1430 \$1462 \$1429 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$96 \$1432 \$1463 \$1431 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$97 \$1371 \$1464 \$1370 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$98 \$1373 \$1465 \$1372 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$99 \$1375 \$1466 \$1374 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$100 \$1377 \$1467 \$1376 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$101 \$1379 \$1468 \$1378 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$102 \$1381 \$1469 \$1380 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$103 \$1383 \$1470 \$1382 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$104 \$1385 \$1471 \$1384 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$105 \$1522 \$1621 \$1521 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$106 \$1524 \$1622 \$1523 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$107 \$1526 \$1623 \$1525 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$108 \$1528 \$1624 \$1527 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$109 \$1530 \$1625 \$1529 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$110 \$1532 \$1626 \$1531 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$111 \$1534 \$1627 \$1533 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$112 \$1536 \$1628 \$1535 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$113 \$1538 \$1629 \$1537 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$114 \$1540 \$1630 \$1539 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$115 \$1542 \$1631 \$1541 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$116 \$1544 \$1632 \$1543 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$117 \$1546 \$1633 \$1545 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$118 \$1548 \$1634 \$1547 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$119 \$1550 \$1635 \$1549 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$120 \$1552 \$1636 \$1551 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$121 \$1554 \$1569 \$1553 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$122 \$1556 \$1570 \$1555 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$123 \$1558 \$1571 \$1557 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$124 \$1560 \$1572 \$1559 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$125 \$1562 \$1573 \$1561 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$126 \$1564 \$1574 \$1563 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$127 \$1566 \$1575 \$1565 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$128 \$1568 \$1576 \$1567 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$129 \$1674 \$1729 \$1673 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$130 \$1676 \$1730 \$1675 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$131 \$1678 \$1731 \$1677 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$132 \$1680 \$1732 \$1679 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$133 \$1682 \$1733 \$1681 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$134 \$1684 \$1734 \$1683 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$135 \$1686 \$1735 \$1685 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$136 \$1688 \$1736 \$1687 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$137 \$1690 \$1737 \$1689 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$138 \$1692 \$1738 \$1691 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$139 \$1694 \$1739 \$1693 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$140 \$1696 \$1740 \$1695 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$141 \$1698 \$1741 \$1697 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$142 \$1700 \$1742 \$1699 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$143 \$1702 \$1743 \$1701 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$144 \$1704 \$1744 \$1703 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$145 \$1643 \$1745 \$1642 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$146 \$1645 \$1746 \$1644 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$147 \$1647 \$1747 \$1646 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$148 \$1649 \$1748 \$1648 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$149 \$1651 \$1749 \$1650 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$150 \$1653 \$1750 \$1652 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$151 \$1655 \$1751 \$1654 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$152 \$1657 \$1752 \$1656 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$153 \$1726 \$1865 \$1725 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$154 \$1728 \$1866 \$1727 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$155 \$1798 \$1867 \$1797 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$156 \$1800 \$1868 \$1799 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$157 \$1802 \$1869 \$1801 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$158 \$1804 \$1870 \$1803 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$159 \$1806 \$1871 \$1805 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$160 \$1808 \$1872 \$1807 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$161 \$1810 \$1873 \$1809 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$162 \$1812 \$1874 \$1811 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$163 \$1814 \$1875 \$1813 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$164 \$1816 \$1876 \$1815 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$165 \$1818 \$1877 \$1817 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$166 \$1820 \$1878 \$1819 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$167 \$1822 \$1879 \$1821 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$168 \$1824 \$1880 \$1823 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$169 \$1826 \$1881 \$1825 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$170 \$1828 \$1882 \$1827 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$171 \$1830 \$1883 \$1829 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$172 \$1832 \$1884 \$1831 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$173 \$1834 \$1885 \$1833 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$174 \$1836 \$1886 \$1835 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$175 \$1838 \$1887 \$1837 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$176 \$1840 \$1888 \$1839 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$177 \$1842 \$1889 \$1841 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$178 \$1844 \$1890 \$1843 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$179 \$1938 \$2009 \$1937 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$180 \$1940 \$2010 \$1939 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$181 \$1942 \$2011 \$1941 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$182 \$1944 \$2012 \$1943 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$183 \$1946 \$2013 \$1945 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$184 \$1948 \$2014 \$1947 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$185 \$1950 \$2015 \$1949 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$186 \$1952 \$2016 \$1951 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$187 \$1954 \$2017 \$1953 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$188 \$1956 \$2018 \$1955 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$189 \$1958 \$2019 \$1957 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$190 \$1960 \$2020 \$1959 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$191 \$1962 \$2021 \$1961 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$192 \$1964 \$2022 \$1963 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$193 \$1966 \$2023 \$1965 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$194 \$1968 \$2024 \$1967 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$195 \$1970 \$2025 \$1969 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$196 \$1972 \$2026 \$1971 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$197 \$1974 \$2027 \$1973 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$198 \$1976 \$2028 \$1975 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$199 \$1978 \$2029 \$1977 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$200 \$1980 \$2030 \$1979 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$201 \$1982 \$2031 \$1981 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$202 \$1984 \$2032 \$1983 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$203 \$1986 \$2033 \$1985 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$204 \$1988 \$2034 \$1987 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$205 \$2118 \$2136 \$2117 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$206 \$2120 \$2137 \$2119 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$207 \$2168 \$2289 \$2167 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$208 \$2170 \$2290 \$2169 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$209 \$2172 \$2291 \$2171 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$210 \$2174 \$2292 \$2173 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$211 \$2191 \$2293 \$2190 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$212 \$2193 \$2294 \$2192 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$213 \$2195 \$2295 \$2194 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$214 \$2197 \$2296 \$2196 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$215 \$2199 \$2297 \$2198 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$216 \$2201 \$2298 \$2200 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$217 \$2203 \$2299 \$2202 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$218 \$2205 \$2300 \$2204 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$219 \$2207 \$2301 \$2206 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$220 \$2209 \$2302 \$2208 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$221 \$2211 \$2303 \$2210 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$222 \$2213 \$2304 \$2212 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$223 \$2215 \$2305 \$2214 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$224 \$2217 \$2306 \$2216 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$225 \$2219 \$2307 \$2218 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$226 \$2221 \$2308 \$2220 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$227 \$2223 \$2309 \$2222 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$228 \$2225 \$2310 \$2224 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$229 \$2087 \$2139 \$2086 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$230 \$2089 \$2140 \$2088 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$231 \$2091 \$2141 \$2090 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$232 \$2093 \$2142 \$2092 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$233 \$2095 \$2143 \$2094 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$234 \$2097 \$2144 \$2096 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$235 \$2099 \$2145 \$2098 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$236 \$2101 \$2146 \$2100 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$237 \$2247 \$2287 \$2246 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$238 \$2249 \$2288 \$2248 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$239 \$2319 \$2425 \$2318 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$240 \$2321 \$2426 \$2320 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$241 \$2323 \$2427 \$2322 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$242 \$2325 \$2428 \$2324 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$243 \$2327 \$2429 \$2326 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$244 \$2329 \$2430 \$2328 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$245 \$2331 \$2431 \$2330 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$246 \$2333 \$2432 \$2332 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$247 \$2335 \$2433 \$2334 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$248 \$2337 \$2434 \$2336 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$249 \$2339 \$2435 \$2338 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$250 \$2341 \$2436 \$2340 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$251 \$2343 \$2437 \$2342 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$252 \$2345 \$2438 \$2344 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$253 \$2347 \$2439 \$2346 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$254 \$2349 \$2440 \$2348 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$255 \$2351 \$2441 \$2350 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$256 \$2353 \$2442 \$2352 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$257 \$2368 \$2443 \$2367 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$258 \$2370 \$2444 \$2369 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$259 \$2372 \$2445 \$2371 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$260 \$2374 \$2446 \$2373 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$261 \$2376 \$2447 \$2375 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$262 \$2378 \$2448 \$2377 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$263 \$2380 \$2449 \$2379 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$264 \$2382 \$2450 \$2381 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$265 \$2384 \$2451 \$2383 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$266 \$2386 \$2452 \$2385 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$267 \$2418 \$2497 \$2417 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$268 \$2420 \$2498 \$2419 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$269 \$2360 \$2421 \$2359 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$270 \$2362 \$2422 \$2361 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$271 \$2364 \$2423 \$2363 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$272 \$2366 \$2424 \$2365 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$273 \$2500 \$2597 \$2499 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$274 \$2502 \$2598 \$2501 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$275 \$2504 \$2599 \$2503 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$276 \$2506 \$2600 \$2505 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$277 \$2508 \$2601 \$2507 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$278 \$2510 \$2602 \$2509 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$279 \$2512 \$2603 \$2511 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$280 \$2514 \$2604 \$2513 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$281 \$2516 \$2605 \$2515 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$282 \$2518 \$2606 \$2517 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$283 \$2520 \$2607 \$2519 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$284 \$2522 \$2608 \$2521 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$285 \$2524 \$2609 \$2523 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$286 \$2526 \$2610 \$2525 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$287 \$2528 \$2611 \$2527 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$288 \$2530 \$2612 \$2529 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$289 \$2532 \$2613 \$2531 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$290 \$2534 \$2614 \$2533 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$291 \$2551 \$2615 \$2550 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$292 \$2553 \$2616 \$2552 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$293 \$2555 \$2617 \$2554 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$294 \$2557 \$2618 \$2556 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$295 \$2559 \$2619 \$2558 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$296 \$2561 \$2620 \$2560 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$297 \$2563 \$2621 \$2562 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$298 \$2565 \$2622 \$2564 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$299 \$2567 \$2623 \$2566 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$300 \$2569 \$2624 \$2568 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$301 \$2586 \$2742 \$2585 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$302 \$2588 \$2743 \$2587 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$303 \$2590 \$2667 \$2589 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$304 \$2592 \$2668 \$2591 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$305 \$2594 \$2669 \$2593 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$306 \$2596 \$2670 \$2595 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$307 \$2672 \$2792 \$2671 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$308 \$2674 \$2793 \$2673 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$309 \$2676 \$2794 \$2675 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$310 \$2678 \$2795 \$2677 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$311 \$2680 \$2796 \$2679 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$312 \$2682 \$2797 \$2681 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$313 \$2684 \$2798 \$2683 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$314 \$2686 \$2799 \$2685 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$315 \$2688 \$2800 \$2687 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$316 \$2690 \$2801 \$2689 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$317 \$2692 \$2802 \$2691 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$318 \$2694 \$2803 \$2693 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$319 \$2696 \$2804 \$2695 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$320 \$2698 \$2805 \$2697 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$321 \$2700 \$2806 \$2699 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$322 \$2702 \$2807 \$2701 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$323 \$2704 \$2808 \$2703 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$324 \$2706 \$2809 \$2705 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$325 \$2708 \$2810 \$2707 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$326 \$2710 \$2811 \$2709 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$327 \$2712 \$2812 \$2711 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$328 \$2714 \$2813 \$2713 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$329 \$2716 \$2814 \$2715 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$330 \$2718 \$2815 \$2717 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$331 \$2720 \$2816 \$2719 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$332 \$2722 \$2817 \$2721 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$333 \$2724 \$2818 \$2723 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$334 \$2726 \$2819 \$2725 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$335 \$2831 \$2890 \$2830 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$336 \$2833 \$2891 \$2832 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$337 \$2785 \$2892 \$2784 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$338 \$2787 \$2893 \$2786 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$339 \$2789 \$2894 \$2788 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$340 \$2791 \$2895 \$2790 \$728 pfet_05v0_dn L=0.5U W=4U AS=3.08P AD=3.08P
+ PS=9.54U PD=9.54U
M$341 \$2840 \$2960 \$2839 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$342 \$2842 \$2961 \$2841 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$343 \$2844 \$2962 \$2843 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$344 \$2846 \$2963 \$2845 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$345 \$2848 \$2964 \$2847 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$346 \$2850 \$2965 \$2849 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$347 \$2852 \$2966 \$2851 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$348 \$2854 \$2967 \$2853 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$349 \$2856 \$2968 \$2855 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$350 \$2858 \$2969 \$2857 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$351 \$2860 \$2970 \$2859 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$352 \$2862 \$2971 \$2861 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$353 \$2864 \$2972 \$2863 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$354 \$2866 \$2973 \$2865 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$355 \$2868 \$2974 \$2867 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$356 \$2870 \$2975 \$2869 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$357 \$2872 \$2976 \$2871 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$358 \$2874 \$2977 \$2873 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$359 \$2897 \$2978 \$2896 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$360 \$2899 \$2979 \$2898 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$361 \$2901 \$2980 \$2900 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$362 \$2903 \$2981 \$2902 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$363 \$2905 \$2982 \$2904 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$364 \$2907 \$2983 \$2906 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$365 \$2909 \$2984 \$2908 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$366 \$2911 \$2985 \$2910 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$367 \$2913 \$2986 \$2912 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$368 \$2915 \$2987 \$2914 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$369 \$3019 \$3159 \$3018 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$370 \$3021 \$3160 \$3020 \$728 pfet_05v0_dn L=3.2U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$371 \$3023 \$3078 \$3022 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$372 \$3025 \$3079 \$3024 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$373 \$3027 \$3080 \$3026 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$374 \$3029 \$3081 \$3028 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$375 \$3031 \$3082 \$3030 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$376 \$3033 \$3083 \$3032 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$377 \$3035 \$3084 \$3034 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$378 \$3037 \$3085 \$3036 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$379 \$3039 \$3086 \$3038 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$380 \$3041 \$3087 \$3040 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$381 \$3043 \$3088 \$3042 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$382 \$3045 \$3089 \$3044 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$383 \$3047 \$3090 \$3046 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$384 \$3049 \$3091 \$3048 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$385 \$3051 \$3092 \$3050 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$386 \$3053 \$3093 \$3052 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$387 \$3055 \$3094 \$3054 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$388 \$3057 \$3095 \$3056 \$728 pfet_05v0_dn L=0.8U W=3.2U AS=2.464P AD=2.464P
+ PS=7.94U PD=7.94U
M$389 \$37 \$45 \$36 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$390 \$39 \$48 \$38 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$391 \$41 \$51 \$40 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$392 \$43 \$54 \$42 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$393 \$46 \$60 \$44 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$394 \$49 \$61 \$47 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$395 \$52 \$62 \$50 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$396 \$55 \$63 \$53 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$397 \$70 \$69 \$68 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$398 \$73 \$72 \$71 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$399 \$76 \$75 \$74 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$400 \$79 \$78 \$77 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P PS=2.46U
+ PD=2.46U
M$401 \$85 \$108 \$84 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$402 \$87 \$109 \$86 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$403 \$89 \$110 \$88 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$404 \$91 \$111 \$90 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$405 \$93 \$112 \$92 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$406 \$95 \$113 \$94 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$407 \$97 \$114 \$96 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$408 \$99 \$115 \$98 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$409 \$101 \$116 \$100 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$410 \$103 \$117 \$102 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$411 \$105 \$118 \$104 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$412 \$107 \$119 \$106 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$413 \$141 \$198 \$140 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$414 \$143 \$199 \$142 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$415 \$145 \$200 \$144 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$416 \$147 \$201 \$146 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$417 \$149 \$202 \$148 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$418 \$151 \$203 \$150 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$419 \$153 \$204 \$152 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$420 \$155 \$205 \$154 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$421 \$157 \$206 \$156 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$422 \$159 \$207 \$158 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$423 \$169 \$222 \$168 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$424 \$171 \$223 \$170 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$425 \$173 \$224 \$172 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$426 \$175 \$225 \$174 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$427 \$177 \$226 \$176 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$428 \$179 \$227 \$178 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$429 \$181 \$228 \$180 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$430 \$183 \$229 \$182 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$431 \$133 \$160 \$132 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$432 \$135 \$161 \$134 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$433 \$137 \$162 \$136 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$434 \$139 \$163 \$138 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$435 \$231 \$292 \$230 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$436 \$233 \$293 \$232 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$437 \$235 \$294 \$234 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$438 \$237 \$295 \$236 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$439 \$239 \$296 \$238 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$440 \$241 \$297 \$240 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$441 \$243 \$298 \$242 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$442 \$245 \$299 \$244 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$443 \$186 \$185 \$184 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$444 \$189 \$188 \$187 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$445 \$192 \$191 \$190 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$446 \$195 \$194 \$193 \$33 nfet_05v0_dn L=2U W=0.5U AS=0.365P AD=0.365P
+ PS=2.46U PD=2.46U
M$447 \$197 \$255 \$196 \$33 nfet_05v0_dn L=4U W=1U AS=0.73P AD=0.73P PS=3.46U
+ PD=3.46U
M$448 \$257 \$318 \$256 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$449 \$259 \$319 \$258 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$450 \$261 \$320 \$260 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$451 \$263 \$321 \$262 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$452 \$265 \$322 \$264 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$453 \$267 \$323 \$266 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$454 \$269 \$324 \$268 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$455 \$271 \$325 \$270 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$456 \$273 \$326 \$272 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$457 \$275 \$327 \$274 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$458 \$277 \$328 \$276 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$459 \$279 \$329 \$278 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$460 \$281 \$330 \$280 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$461 \$283 \$331 \$282 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$462 \$285 \$332 \$284 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$463 \$287 \$333 \$286 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$464 \$289 \$334 \$288 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$465 \$291 \$335 \$290 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$466 \$337 \$396 \$336 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$467 \$339 \$397 \$338 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$468 \$341 \$398 \$340 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$469 \$343 \$399 \$342 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$470 \$345 \$400 \$344 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$471 \$347 \$401 \$346 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$472 \$349 \$402 \$348 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$473 \$351 \$403 \$350 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$474 \$361 \$412 \$360 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$475 \$363 \$413 \$362 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$476 \$365 \$414 \$364 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$477 \$367 \$415 \$366 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$478 \$369 \$416 \$368 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$479 \$371 \$417 \$370 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$480 \$373 \$418 \$372 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$481 \$375 \$419 \$374 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$482 \$377 \$420 \$376 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$483 \$379 \$421 \$378 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$484 \$381 \$432 \$380 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$485 \$383 \$433 \$382 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$486 \$385 \$434 \$384 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$487 \$387 \$435 \$386 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$488 \$389 \$436 \$388 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$489 \$391 \$437 \$390 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$490 \$393 \$438 \$392 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$491 \$395 \$439 \$394 \$33 nfet_05v0_dn L=1U W=4U AS=2.92P AD=2.92P PS=9.46U
+ PD=9.46U
M$492 \$441 \$484 \$440 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$493 \$443 \$485 \$442 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$494 \$445 \$486 \$444 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$495 \$447 \$487 \$446 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$496 \$449 \$488 \$448 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$497 \$451 \$489 \$450 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$498 \$453 \$490 \$452 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$499 \$455 \$491 \$454 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$500 \$465 \$526 \$464 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$501 \$467 \$527 \$466 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$502 \$469 \$528 \$468 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$503 \$471 \$529 \$470 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$504 \$473 \$530 \$472 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$505 \$475 \$531 \$474 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$506 \$477 \$532 \$476 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$507 \$479 \$533 \$478 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$508 \$481 \$534 \$480 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$509 \$483 \$535 \$482 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$510 \$511 \$556 \$510 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$511 \$513 \$557 \$512 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$512 \$515 \$558 \$514 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$513 \$517 \$559 \$516 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$514 \$519 \$560 \$518 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$515 \$521 \$561 \$520 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$516 \$523 \$562 \$522 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$517 \$525 \$563 \$524 \$33 nfet_05v0_dn L=1U W=3.2U AS=2.336P AD=2.336P
+ PS=7.86U PD=7.86U
M$518 \$537 \$614 \$536 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$519 \$539 \$615 \$538 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$520 \$541 \$616 \$540 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$521 \$543 \$617 \$542 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$522 \$545 \$618 \$544 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$523 \$547 \$619 \$546 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$524 \$549 \$620 \$548 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$525 \$551 \$621 \$550 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$526 \$553 \$622 \$552 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$527 \$555 \$623 \$554 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$528 \$633 \$652 \$632 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$529 \$635 \$653 \$634 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$530 \$637 \$654 \$636 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$531 \$639 \$655 \$638 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$532 \$641 \$656 \$640 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$533 \$643 \$657 \$642 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$534 \$645 \$658 \$644 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$535 \$647 \$659 \$646 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$536 \$649 \$660 \$648 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
M$537 \$651 \$661 \$650 \$33 nfet_05v0_dn L=0.6U W=4U AS=2.92P AD=2.92P
+ PS=9.46U PD=9.46U
Q$538 I1_default_C I1_default_B I1_default_E pnp_05p00x05p00 AE=1200P PE=960U
+ AB=41.9904P PB=25.92U AC=41.9904P PC=25.92U NE=48
R$586 \$4 \$5 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$587 \$7 \$8 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$588 \$10 \$11 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$589 \$13 \$14 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$590 \$18 \$19 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$591 \$21 \$22 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$592 \$26 \$27 SUB 4500 ppolyf_u_1k L=4.5U W=1U
R$593 \$29 \$30 SUB 4500 ppolyf_u_1k L=4.5U W=1U
.ENDS bandgap
