* NGSPICE file created from test_decoder.ext - technology: gf180mcuD

.subckt test_decoder VDD VSS EN SEL[0] SEL[1] SEL[2] EN0 EN1 EN2 EN3 EN4 EN5 EN6 EN7
X0 VSS a_n56986_5965# a_n56986_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X1 VDD a_n47266_6815# a_n47266_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X2 VDD SEL[1] a_n44836_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X3 VDD a_n47266_3415# a_n47266_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X4 VDD a_n49696_5115# a_n49696_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X5 VSS a_n52126_5115# a_n52126_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X6 VDD a_n39976_5115# a_n39976_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X7 VSS EN a_n49696_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X8 VDD EN a_n54556_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X9 a_n56986_8515# a_n56986_6815# a_n56986_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X10 VDD a_n42406_6815# a_n42406_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X11 VSS a_n54556_5115# a_n54556_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X12 VSS EN a_n44836_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X13 VDD SEL[2] a_n42406_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X14 a_n52126_8515# a_n52126_6815# a_n52126_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X15 VDD a_n44836_5115# a_n44836_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X16 VSS a_n39976_5115# a_n39976_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X17 VDD SEL[1] a_n49696_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X18 VSS EN a_n47266_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X19 VSS a_n49696_7665# EN3 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X20 VDD SEL[1] a_n39976_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X21 a_n54556_8515# a_n54556_6815# a_n54556_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X22 VSS EN a_n42406_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X23 VSS a_n44836_7665# EN5 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X24 VDD SEL[1] a_n47266_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X25 VDD a_n56986_6815# a_n56986_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X26 VDD a_n56986_3415# a_n56986_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X27 a_n39976_8515# a_n39976_6815# a_n39976_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X28 VDD a_n44836_1715# a_n44836_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X29 VSS a_n47266_7665# EN4 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X30 VSS a_n42406_7665# EN6 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X31 VDD SEL[0] a_n42406_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X32 VDD a_n47266_5115# a_n47266_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X33 VDD a_n52126_6815# a_n52126_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X34 VDD a_n52126_2565# a_n52126_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X35 VSS a_n49696_5115# a_n49696_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X36 VSS SEL[2] a_n56986_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X37 VSS a_n56986_4265# a_n56986_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X38 VSS a_n44836_5115# a_n44836_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X39 VDD a_n42406_5115# a_n42406_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X40 VDD SEL[0] a_n56986_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X41 a_n52126_5965# a_n52126_4265# a_n52126_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X42 VSS a_n51980_5905# a_n52126_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X43 VDD a_n47266_1715# a_n47266_3415# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X44 VDD SEL[2] a_n49696_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X45 a_n49696_8515# a_n49696_6815# a_n49696_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X46 VDD SEL[2] a_n39976_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X47 VSS a_n47266_5115# a_n47266_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X48 a_n44836_8515# a_n44836_6815# a_n44836_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X49 VDD a_n54556_6815# a_n54556_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X50 a_n54556_5965# a_n54556_4265# a_n54556_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X51 VSS SEL[2] a_n54556_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X52 VSS a_n42406_5115# a_n42406_6815# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X53 VDD SEL[0] a_n52126_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X54 VDD a_n54556_3415# a_n54556_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X55 VDD a_n56986_5965# a_n56986_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X56 VDD a_n42406_1715# a_n42406_3415# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X57 VSS SEL[2] a_n39976_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X58 VDD SEL[2] a_n44836_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X59 a_n39976_5965# a_n39976_4265# a_n39976_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X60 a_n47266_8515# a_n47266_6815# a_n47266_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X61 a_n42406_8515# a_n42406_6815# a_n42406_7665# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X62 VDD a_n52126_5115# a_n52126_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X63 VDD a_n56986_1715# a_n56986_3415# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X64 VSS a_n56986_1715# a_n56986_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X65 VDD SEL[0] a_n54556_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X66 VDD a_n47266_4265# a_n47266_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X67 VSS SEL[1] a_n52126_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X68 VDD SEL[1] a_n52126_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X69 a_n49696_5965# a_n49696_4265# a_n49696_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X70 VSS SEL[2] a_n49696_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X71 a_n56986_5115# a_n56986_3415# a_n56986_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X72 a_n44836_5965# a_n44836_4265# a_n44836_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X73 VSS SEL[2] a_n44836_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X74 VDD a_n54556_5115# a_n54556_6815# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X75 VSS a_n54556_1715# a_n54556_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X76 VSS a_n52126_2565# a_n52126_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X77 VDD a_n42406_4265# a_n42406_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X78 VSS SEL[1] a_n39976_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X79 VDD a_n49696_4265# a_n49696_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X80 a_n47266_5965# SEL[0] a_n47266_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X81 VSS a_n47266_4265# a_n47266_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X82 VDD a_n39976_4265# a_n39976_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X83 VSS a_n54556_3415# a_n54556_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X84 a_n42406_5965# a_n42406_3415# a_n42406_5115# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X85 VSS a_n42406_4265# a_n42406_5965# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X86 VDD a_n54556_1715# a_n54556_3415# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X87 VDD a_n56986_4265# a_n56986_5965# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X88 VSS a_n39976_2565# a_n39976_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X89 VDD a_n49696_7665# EN3 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X90 VDD a_n39976_7665# EN7 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X91 VDD a_n44836_4265# a_n44836_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X92 a_n56986_2565# SEL[0] a_n56986_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X93 VSS SEL[0] a_n52126_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X94 VDD a_n44836_7665# EN5 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X95 VDD a_n51980_5905# a_n52126_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X96 VDD a_n49696_1715# a_n49696_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X97 VSS SEL[1] a_n49696_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X98 VDD SEL[0] a_n39976_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X99 a_n54556_2565# SEL[0] a_n54556_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X100 VSS SEL[1] a_n56986_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X101 VSS a_n44836_1715# a_n44836_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X102 a_n52126_3415# a_n52126_1715# a_n52126_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X103 VSS SEL[2] a_n51980_5905# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X104 VDD SEL[0] a_n44836_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X105 VDD SEL[0] a_n47266_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X106 VSS a_n49696_2565# a_n49696_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X107 VSS a_n47266_1715# a_n47266_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X108 VSS SEL[1] a_n54556_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X109 VSS a_n42406_1715# a_n42406_3415# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X110 VSS a_n44836_2565# a_n44836_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X111 VDD a_n47266_7665# EN4 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X112 VDD SEL[2] a_n54556_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X113 a_n39976_3415# SEL[0] a_n39976_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X114 VDD a_n42406_3415# a_n42406_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X115 VSS a_n47266_3415# a_n47266_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X116 VSS SEL[2] a_n42406_4265# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X117 VDD a_n42406_7665# EN6 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X118 VDD SEL[2] a_n47266_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X119 VDD EN a_n49696_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X120 VDD SEL[2] a_n56986_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X121 VSS SEL[0] a_n49696_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X122 VDD EN a_n39976_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X123 VSS SEL[1] a_n44836_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X124 VDD a_n56986_7665# EN0 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X125 VDD SEL[1] a_n42406_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X126 VDD EN a_n44836_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X127 VDD a_n52126_4265# a_n52126_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X128 a_n47266_2565# SEL[1] a_n47266_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X129 a_n49696_3415# a_n49696_1715# a_n49696_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X130 a_n42406_2565# SEL[0] a_n42406_1715# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X131 a_n44836_3415# SEL[0] a_n44836_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X132 VDD a_n52126_7665# EN2 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X133 VDD SEL[1] a_n56986_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X134 VSS SEL[2] a_n47266_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X135 VSS SEL[1] a_n42406_2565# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X136 VDD a_n54556_4265# a_n54556_5115# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X137 VDD EN a_n47266_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X138 VDD a_n52126_1715# a_n52126_2565# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X139 VDD a_n54556_7665# EN1 VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X140 VDD EN a_n42406_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X141 VSS EN a_n56986_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X142 VDD a_n49696_6815# a_n49696_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X143 VDD a_n49696_2565# a_n49696_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X144 VSS EN a_n52126_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X145 VDD a_n39976_2565# a_n39976_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X146 VDD a_n39976_6815# a_n39976_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X147 VDD SEL[1] a_n54556_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X148 VSS EN a_n54556_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X149 VSS a_n56986_7665# EN0 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X150 VDD EN a_n56986_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X151 VDD a_n44836_2565# a_n44836_4265# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X152 VDD a_n44836_6815# a_n44836_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X153 VSS a_n52126_7665# EN2 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X154 VSS EN a_n39976_8515# VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X155 VSS a_n54556_7665# EN1 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
X156 VDD EN a_n52126_7665# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X157 VDD SEL[0] a_n49696_1715# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X158 VDD SEL[2] a_n51980_5905# VDD pfet_05v0 ad=0.385p pd=2.54u as=0.385p ps=2.54u w=0.5u l=0.5u
X159 VSS a_n39976_7665# EN7 VSS nfet_05v0 ad=0.365p pd=2.46u as=0.365p ps=2.46u w=0.5u l=0.6u
.ends

