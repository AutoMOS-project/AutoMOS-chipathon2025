* Extracted by KLayout with GF180MCU LVS runset on : 12/09/2025 06:22

.SUBCKT ldo VSS VDD VOUT IBIAS LDO_EN VFB VREF
M$1 VDD LDO_EN \$506 VDD pfet_05v0_dn L=0.5U W=0.6U AS=0.462P AD=0.462P
+ PS=2.74U PD=2.74U
M$2 VDD \$506 \$182 VDD pfet_05v0_dn L=0.5U W=0.6U AS=0.462P AD=0.462P PS=2.74U
+ PD=2.74U
M$3 VDD \$182 \$2652 VDD pfet_05v0_dn L=0.5U W=2U AS=1.54P AD=1.54P PS=5.54U
+ PD=5.54U
M$4 VDD \$182 \$2128 VDD pfet_05v0_dn L=0.5U W=2U AS=1.54P AD=1.54P PS=5.54U
+ PD=5.54U
M$5 VDD \$182 \$181 VDD pfet_05v0_dn L=0.5U W=2U AS=1.54P AD=1.54P PS=5.54U
+ PD=5.54U
M$6 VDD \$181 VOUT VDD pfet_05v0_dn L=0.5U W=500U AS=385P AD=385P PS=1015.4U
+ PD=1015.4U
M$16 VDD VDD VDD VDD pfet_05v0_dn L=1U W=110U AS=84.7P AD=84.7P PS=250.8U
+ PD=250.8U
M$18 VDD \$2652 \$181 VDD pfet_05v0_dn L=1U W=33U AS=25.41P AD=25.41P PS=75.24U
+ PD=75.24U
M$23 VDD \$2128 \$2128 VDD pfet_05v0_dn L=1U W=11U AS=8.47P AD=8.47P PS=25.08U
+ PD=25.08U
M$24 VDD \$2128 \$42 VDD pfet_05v0_dn L=1U W=11U AS=8.47P AD=8.47P PS=25.08U
+ PD=25.08U
M$27 VDD \$2652 \$2652 VDD pfet_05v0_dn L=1U W=11U AS=8.47P AD=8.47P PS=25.08U
+ PD=25.08U
M$48 VSS VSS VSS VSS nfet_05v0_dn L=1U W=56U AS=40.88P AD=40.88P PS=152.88U
+ PD=152.88U
M$55 VSS \$42 \$181 VSS nfet_05v0_dn L=1U W=7.5U AS=5.475P AD=5.475P PS=23.76U
+ PD=23.76U
M$57 VSS \$42 \$42 VSS nfet_05v0_dn L=1U W=2.5U AS=1.825P AD=1.825P PS=7.92U
+ PD=7.92U
M$74 VSS \$125 \$114 VSS nfet_05v0_dn L=1U W=6U AS=4.38P AD=4.38P PS=14.92U
+ PD=14.92U
M$77 VSS \$125 \$125 VSS nfet_05v0_dn L=1U W=6U AS=4.38P AD=4.38P PS=14.92U
+ PD=14.92U
M$88 VSS \$506 \$42 VSS nfet_05v0_dn L=0.6U W=2U AS=1.46P AD=1.46P PS=5.46U
+ PD=5.46U
M$89 VSS \$506 \$125 VSS nfet_05v0_dn L=0.6U W=2U AS=1.46P AD=1.46P PS=5.46U
+ PD=5.46U
M$90 \$125 \$182 IBIAS VSS nfet_05v0_dn L=0.6U W=2U AS=1.46P AD=1.46P PS=5.46U
+ PD=5.46U
M$91 VSS VSS VSS VSS nfet_05v0_dn L=0.6U W=130U AS=94.9P AD=94.9P PS=297.96U
+ PD=297.96U
M$92 VSS LDO_EN \$506 VSS nfet_05v0_dn L=0.6U W=0.42U AS=0.315P AD=0.315P
+ PS=2.34U PD=2.34U
M$93 VSS \$506 \$182 VSS nfet_05v0_dn L=0.6U W=0.42U AS=0.315P AD=0.315P
+ PS=2.34U PD=2.34U
M$103 \$114 VREF \$2128 VSS nfet_05v0_dn L=0.6U W=70U AS=51.1P AD=51.1P
+ PS=160.44U PD=160.44U
M$104 \$114 VFB \$2652 VSS nfet_05v0_dn L=0.6U W=70U AS=51.1P AD=51.1P
+ PS=160.44U PD=160.44U
C$147 \$179 \$181 5e-12 cap_mim_2f0_m4m5_noshield A=2500P P=400U
.ENDS ldo
