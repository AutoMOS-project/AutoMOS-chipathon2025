** sch_path: /home/vasil/Downloads/AutoMOS-chipathon2025/designs/Chipathon2025_pads/xschem/io_secondary_AC_tb.sch
**.subckt io_secondary_AC_tb
V1 DVDD GND 5
V2 VDD GND 5
V3 DVSS GND 0
V4 VSS GND 0
V5 net1 GND DC 3 AC 1
R1 PAD net1 1k m=1
XIO1 DVSS DVDD VSS VDD PAD asig gf180mcu_fd_io__asig_5p0_extracted
XIO2 VDD to_gate asig VSS io_secondary_5p0
**** begin user architecture code

.include /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice diode_typical
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical



.control
   save all
   ac dec 100 1k 100G

   write io_secondary_AC.raw
* run
* display
* plot PAD ASIG
* plot vdb(asig) vdb(to_gate)
.endc



.include /home/vasil/Downloads/AutoMOS-chipathon2025/designs/Chipathon2025_pads/xschem/gf180mcu_fd_io__asig_5p0_extracted.spice

**** end user architecture code
**.ends

* expanding   symbol:  Chipathon2025_pads/xschem/symbols/io_secondary_5p0/io_secondary_5p0.sym # of pins=4
** sym_path: /home/vasil/Downloads/AutoMOS-chipathon2025/designs/Chipathon2025_pads/xschem/symbols/io_secondary_5p0/io_secondary_5p0.sym
** sch_path: /home/vasil/Downloads/AutoMOS-chipathon2025/designs/Chipathon2025_pads/xschem/symbols/io_secondary_5p0/io_secondary_5p0.sch
.subckt io_secondary_5p0 VDD to_gate ASIG5V VSS


*.iopin VSS
*.iopin VDD
*.iopin to_gate
*.iopin ASIG5V
D1 to_gate VDD diode_pd2nw_06v0 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
XR1 to_gate ASIG5V VDD ppolyf_u r_width=16e-6 r_length=4e-6 m=1
D2 VSS to_gate diode_nd2ps_06v0 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
.ends

.GLOBAL GND
.end
